module rom_1p #(
	int Depth, 
 	int DATA_WIDTH = 32, 
 	int ADDR_WIDTH = 32 
 ) (
	input logic clk_i, 
	input logic req_i, 
	input logic [ADDR_WIDTH-1:0] addr_i, 
	output logic [DATA_WIDTH-1:0] data_o 
 );
	always_ff @(posedge clk_i) begin
		case (addr_i)
			32'h00100000 : data_o = 32'h0eb0006f ;
			32'h00100004 : data_o = 32'h0e70006f ;
			32'h00100008 : data_o = 32'h0e30006f ;
			32'h0010000c : data_o = 32'h0df0006f ;
			32'h00100010 : data_o = 32'h0db0006f ;
			32'h00100014 : data_o = 32'h0d70006f ;
			32'h00100018 : data_o = 32'h0d30006f ;
			32'h0010001c : data_o = 32'h0cf0006f ;
			32'h00100020 : data_o = 32'h0cb0006f ;
			32'h00100024 : data_o = 32'h0c70006f ;
			32'h00100028 : data_o = 32'h0c30006f ;
			32'h0010002c : data_o = 32'h0bf0006f ;
			32'h00100030 : data_o = 32'h0bb0006f ;
			32'h00100034 : data_o = 32'h0b70006f ;
			32'h00100038 : data_o = 32'h0b30006f ;
			32'h0010003c : data_o = 32'h0af0006f ;
			32'h00100040 : data_o = 32'h0ab0006f ;
			32'h00100044 : data_o = 32'h0400006f ;
			32'h00100048 : data_o = 32'h0a30006f ;
			32'h0010004c : data_o = 32'h09f0006f ;
			32'h00100050 : data_o = 32'h09b0006f ;
			32'h00100054 : data_o = 32'h0970006f ;
			32'h00100058 : data_o = 32'h0930006f ;
			32'h0010005c : data_o = 32'h08f0006f ;
			32'h00100060 : data_o = 32'h08b0006f ;
			32'h00100064 : data_o = 32'h0870006f ;
			32'h00100068 : data_o = 32'h0830006f ;
			32'h0010006c : data_o = 32'h07f0006f ;
			32'h00100070 : data_o = 32'h07b0006f ;
			32'h00100074 : data_o = 32'h0770006f ;
			32'h00100078 : data_o = 32'h0730006f ;
			32'h0010007c : data_o = 32'h06f0006f ;
			32'h00100080 : data_o = 32'h6410006f ;
			32'h00100084 : data_o = 32'hc686715d ;
			32'h00100088 : data_o = 32'hc29ac496 ;
			32'h0010008c : data_o = 32'hde22c09e ;
			32'h00100090 : data_o = 32'hda2edc2a ;
			32'h00100094 : data_o = 32'hd636d832 ;
			32'h00100098 : data_o = 32'hd23ed43a ;
			32'h0010009c : data_o = 32'hce46d042 ;
			32'h001000a0 : data_o = 32'hca76cc72 ;
			32'h001000a4 : data_o = 32'hc67ec87a ;
			32'h001000a8 : data_o = 32'h00ef0880 ;
			32'h001000ac : data_o = 32'h872a5130 ;
			32'h001000b0 : data_o = 32'h00100797 ;
			32'h001000b4 : data_o = 32'hf6478793 ;
			32'h001000b8 : data_o = 32'h0797c398 ;
			32'h001000bc : data_o = 32'h87930010 ;
			32'h001000c0 : data_o = 32'h4705f5e7 ;
			32'h001000c4 : data_o = 32'h0001c398 ;
			32'h001000c8 : data_o = 32'h42a640b6 ;
			32'h001000cc : data_o = 32'h43864316 ;
			32'h001000d0 : data_o = 32'h55625472 ;
			32'h001000d4 : data_o = 32'h564255d2 ;
			32'h001000d8 : data_o = 32'h572256b2 ;
			32'h001000dc : data_o = 32'h58025792 ;
			32'h001000e0 : data_o = 32'h4e6248f2 ;
			32'h001000e4 : data_o = 32'h4f424ed2 ;
			32'h001000e8 : data_o = 32'h61614fb2 ;
			32'h001000ec : data_o = 32'h30200073 ;
			32'h001000f0 : data_o = 32'hd6067179 ;
			32'h001000f4 : data_o = 32'h1800d422 ;
			32'h001000f8 : data_o = 32'hfca42e23 ;
			32'h001000fc : data_o = 32'hfe042623 ;
			32'h00100100 : data_o = 32'h2783a839 ;
			32'h00100104 : data_o = 32'h2703fec4 ;
			32'h00100108 : data_o = 32'h97bafdc4 ;
			32'h0010010c : data_o = 32'h0007c783 ;
			32'h00100110 : data_o = 32'h2b3d853e ;
			32'h00100114 : data_o = 32'hfec42783 ;
			32'h00100118 : data_o = 32'h26230785 ;
			32'h0010011c : data_o = 32'h2783fef4 ;
			32'h00100120 : data_o = 32'h2703fec4 ;
			32'h00100124 : data_o = 32'h97bafdc4 ;
			32'h00100128 : data_o = 32'h0007c783 ;
			32'h0010012c : data_o = 32'h0001fbf9 ;
			32'h00100130 : data_o = 32'h50b20001 ;
			32'h00100134 : data_o = 32'h61455422 ;
			32'h00100138 : data_o = 32'h71798082 ;
			32'h0010013c : data_o = 32'hd422d606 ;
			32'h00100140 : data_o = 32'h832a1800 ;
			32'h00100144 : data_o = 32'h853288ae ;
			32'h00100148 : data_o = 32'h863a85b6 ;
			32'h0010014c : data_o = 32'h874286be ;
			32'h00100150 : data_o = 32'h0fa3879a ;
			32'h00100154 : data_o = 32'h87c6fcf4 ;
			32'h00100158 : data_o = 32'hfcf40f23 ;
			32'h0010015c : data_o = 32'h0ea387aa ;
			32'h00100160 : data_o = 32'h87aefcf4 ;
			32'h00100164 : data_o = 32'hfcf40e23 ;
			32'h00100168 : data_o = 32'h0da387b2 ;
			32'h0010016c : data_o = 32'h87b6fcf4 ;
			32'h00100170 : data_o = 32'hfcf40d23 ;
			32'h00100174 : data_o = 32'h0ca387ba ;
			32'h00100178 : data_o = 32'h4505fcf4 ;
			32'h0010017c : data_o = 32'h4ab000ef ;
			32'h00100180 : data_o = 32'hfdf44783 ;
			32'h00100184 : data_o = 32'h01879713 ;
			32'h00100188 : data_o = 32'hfde44783 ;
			32'h0010018c : data_o = 32'h8f5d07c2 ;
			32'h00100190 : data_o = 32'hfdd44783 ;
			32'h00100194 : data_o = 32'h8f5d07a2 ;
			32'h00100198 : data_o = 32'hfdc44783 ;
			32'h0010019c : data_o = 32'h26238fd9 ;
			32'h001001a0 : data_o = 32'h4505fef4 ;
			32'h001001a4 : data_o = 32'h4a1000ef ;
			32'h001001a8 : data_o = 32'hfd944683 ;
			32'h001001ac : data_o = 32'hfda44703 ;
			32'h001001b0 : data_o = 32'hfdb44783 ;
			32'h001001b4 : data_o = 32'h85be863a ;
			32'h001001b8 : data_o = 32'hfec42503 ;
			32'h001001bc : data_o = 32'h4a9000ef ;
			32'h001001c0 : data_o = 32'h50b20001 ;
			32'h001001c4 : data_o = 32'h61455422 ;
			32'h001001c8 : data_o = 32'h11018082 ;
			32'h001001cc : data_o = 32'hcc22ce06 ;
			32'h001001d0 : data_o = 32'h8eaa1000 ;
			32'h001001d4 : data_o = 32'h83328e2e ;
			32'h001001d8 : data_o = 32'h85ba8536 ;
			32'h001001dc : data_o = 32'h86c2863e ;
			32'h001001e0 : data_o = 32'h87f68746 ;
			32'h001001e4 : data_o = 32'hfef407a3 ;
			32'h001001e8 : data_o = 32'h072387f2 ;
			32'h001001ec : data_o = 32'h879afef4 ;
			32'h001001f0 : data_o = 32'hfef406a3 ;
			32'h001001f4 : data_o = 32'h062387aa ;
			32'h001001f8 : data_o = 32'h87aefef4 ;
			32'h001001fc : data_o = 32'hfef405a3 ;
			32'h00100200 : data_o = 32'h052387b2 ;
			32'h00100204 : data_o = 32'h87b6fef4 ;
			32'h00100208 : data_o = 32'hfef404a3 ;
			32'h0010020c : data_o = 32'h042387ba ;
			32'h00100210 : data_o = 32'h4505fef4 ;
			32'h00100214 : data_o = 32'h2a5000ef ;
			32'h00100218 : data_o = 32'hfec44683 ;
			32'h0010021c : data_o = 32'hfed44603 ;
			32'h00100220 : data_o = 32'hfee44703 ;
			32'h00100224 : data_o = 32'hfef44783 ;
			32'h00100228 : data_o = 32'h853e85ba ;
			32'h0010022c : data_o = 32'h2ab000ef ;
			32'h00100230 : data_o = 32'hfe844683 ;
			32'h00100234 : data_o = 32'hfe944603 ;
			32'h00100238 : data_o = 32'hfea44703 ;
			32'h0010023c : data_o = 32'hfeb44783 ;
			32'h00100240 : data_o = 32'h853e85ba ;
			32'h00100244 : data_o = 32'h2e9000ef ;
			32'h00100248 : data_o = 32'h853e401c ;
			32'h0010024c : data_o = 32'h337000ef ;
			32'h00100250 : data_o = 32'h353000ef ;
			32'h00100254 : data_o = 32'he789401c ;
			32'h00100258 : data_o = 32'h365000ef ;
			32'h0010025c : data_o = 32'ha00d87aa ;
			32'h00100260 : data_o = 32'h47894018 ;
			32'h00100264 : data_o = 32'h00f71663 ;
			32'h00100268 : data_o = 32'h36d000ef ;
			32'h0010026c : data_o = 32'ha80987aa ;
			32'h00100270 : data_o = 32'h47854018 ;
			32'h00100274 : data_o = 32'h00f71663 ;
			32'h00100278 : data_o = 32'h375000ef ;
			32'h0010027c : data_o = 32'ha00987aa ;
			32'h00100280 : data_o = 32'h40f2853e ;
			32'h00100284 : data_o = 32'h61054462 ;
			32'h00100288 : data_o = 32'h71798082 ;
			32'h0010028c : data_o = 32'hd422d606 ;
			32'h00100290 : data_o = 32'h87aa1800 ;
			32'h00100294 : data_o = 32'h873286ae ;
			32'h00100298 : data_o = 32'hfcf40fa3 ;
			32'h0010029c : data_o = 32'h0f2387b6 ;
			32'h001002a0 : data_o = 32'h87bafcf4 ;
			32'h001002a4 : data_o = 32'hfcf40ea3 ;
			32'h001002a8 : data_o = 32'hfdf44783 ;
			32'h001002ac : data_o = 32'hf713078e ;
			32'h001002b0 : data_o = 32'h47830187 ;
			32'h001002b4 : data_o = 32'h0796fde4 ;
			32'h001002b8 : data_o = 32'h47838f5d ;
			32'h001002bc : data_o = 32'h078afdd4 ;
			32'h001002c0 : data_o = 32'h8fd98b91 ;
			32'h001002c4 : data_o = 32'hfef42623 ;
			32'h001002c8 : data_o = 32'hfec42503 ;
			32'h001002cc : data_o = 32'h339000ef ;
			32'h001002d0 : data_o = 32'h853e87aa ;
			32'h001002d4 : data_o = 32'h542250b2 ;
			32'h001002d8 : data_o = 32'h80826145 ;
			32'h001002dc : data_o = 32'hd6067179 ;
			32'h001002e0 : data_o = 32'h1800d422 ;
			32'h001002e4 : data_o = 32'hfca42e23 ;
			32'h001002e8 : data_o = 32'hfdc42783 ;
			32'h001002ec : data_o = 32'hfef42423 ;
			32'h001002f0 : data_o = 32'hfe042623 ;
			32'h001002f4 : data_o = 32'h2703a835 ;
			32'h001002f8 : data_o = 32'h47a9fe84 ;
			32'h001002fc : data_o = 32'h02f777b3 ;
			32'h00100300 : data_o = 32'h0ff7f793 ;
			32'h00100304 : data_o = 32'h03078793 ;
			32'h00100308 : data_o = 32'h0ff7f713 ;
			32'h0010030c : data_o = 32'hfec42783 ;
			32'h00100310 : data_o = 32'h97a217c1 ;
			32'h00100314 : data_o = 32'hfee78a23 ;
			32'h00100318 : data_o = 32'hfe842703 ;
			32'h0010031c : data_o = 32'h57b347a9 ;
			32'h00100320 : data_o = 32'h242302f7 ;
			32'h00100324 : data_o = 32'h2783fef4 ;
			32'h00100328 : data_o = 32'h0785fec4 ;
			32'h0010032c : data_o = 32'hfef42623 ;
			32'h00100330 : data_o = 32'hfec42703 ;
			32'h00100334 : data_o = 32'hd0e3478d ;
			32'h00100338 : data_o = 32'h478dfce7 ;
			32'h0010033c : data_o = 32'hfef42623 ;
			32'h00100340 : data_o = 32'h2783a831 ;
			32'h00100344 : data_o = 32'h17c1fec4 ;
			32'h00100348 : data_o = 32'hc78397a2 ;
			32'h0010034c : data_o = 32'h853eff47 ;
			32'h00100350 : data_o = 32'h27832601 ;
			32'h00100354 : data_o = 32'h17fdfec4 ;
			32'h00100358 : data_o = 32'hfef42623 ;
			32'h0010035c : data_o = 32'hfec42783 ;
			32'h00100360 : data_o = 32'hfe07d1e3 ;
			32'h00100364 : data_o = 32'h00010001 ;
			32'h00100368 : data_o = 32'h542250b2 ;
			32'h0010036c : data_o = 32'h80826145 ;
			32'h00100370 : data_o = 32'hde067139 ;
			32'h00100374 : data_o = 32'h0080dc22 ;
			32'h00100378 : data_o = 32'h911672f9 ;
			32'h0010037c : data_o = 32'h17c177f9 ;
			32'h00100380 : data_o = 32'h171797a2 ;
			32'h00100384 : data_o = 32'h07130000 ;
			32'h00100388 : data_o = 32'h17b1d067 ;
			32'h0010038c : data_o = 32'h670986ba ;
			32'h00100390 : data_o = 32'h85b6863a ;
			32'h00100394 : data_o = 32'h00ef853e ;
			32'h00100398 : data_o = 32'h07a33ab0 ;
			32'h0010039c : data_o = 32'h47b1fe04 ;
			32'h001003a0 : data_o = 32'hfef40723 ;
			32'h001003a4 : data_o = 32'h06a347e1 ;
			32'h001003a8 : data_o = 32'h0793fef4 ;
			32'h001003ac : data_o = 32'h06230220 ;
			32'h001003b0 : data_o = 32'h05a3fef4 ;
			32'h001003b4 : data_o = 32'h0523fe04 ;
			32'h001003b8 : data_o = 32'h04a3fe04 ;
			32'h001003bc : data_o = 32'h0423fe04 ;
			32'h001003c0 : data_o = 32'h03a3fe04 ;
			32'h001003c4 : data_o = 32'h4803fe04 ;
			32'h001003c8 : data_o = 32'h4783fe74 ;
			32'h001003cc : data_o = 32'h4703fe84 ;
			32'h001003d0 : data_o = 32'h4683feb4 ;
			32'h001003d4 : data_o = 32'h4603fec4 ;
			32'h001003d8 : data_o = 32'h4583fed4 ;
			32'h001003dc : data_o = 32'h4503fee4 ;
			32'h001003e0 : data_o = 32'h3ba1fef4 ;
			32'h001003e4 : data_o = 32'hfe744683 ;
			32'h001003e8 : data_o = 32'hfe844703 ;
			32'h001003ec : data_o = 32'hfeb44783 ;
			32'h001003f0 : data_o = 32'h85ba8636 ;
			32'h001003f4 : data_o = 32'h3d51853e ;
			32'h001003f8 : data_o = 32'hfea42023 ;
			32'h001003fc : data_o = 32'h2c894529 ;
			32'h00100400 : data_o = 32'h2a114501 ;
			32'h00100404 : data_o = 32'h17c177f9 ;
			32'h00100408 : data_o = 32'ha42397a2 ;
			32'h0010040c : data_o = 32'h77f9fe07 ;
			32'h00100410 : data_o = 32'h97a217c1 ;
			32'h00100414 : data_o = 32'hfe87c503 ;
			32'h00100418 : data_o = 32'h17c177f9 ;
			32'h0010041c : data_o = 32'hc58397a2 ;
			32'h00100420 : data_o = 32'h77f9fe87 ;
			32'h00100424 : data_o = 32'h97a217c1 ;
			32'h00100428 : data_o = 32'hfe87c603 ;
			32'h0010042c : data_o = 32'h17c177f9 ;
			32'h00100430 : data_o = 32'hc68397a2 ;
			32'h00100434 : data_o = 32'h77f9fe87 ;
			32'h00100438 : data_o = 32'h97a217c1 ;
			32'h0010043c : data_o = 32'hfe87c703 ;
			32'h00100440 : data_o = 32'h17c177f9 ;
			32'h00100444 : data_o = 32'hc30397a2 ;
			32'h00100448 : data_o = 32'h77f9fe87 ;
			32'h0010044c : data_o = 32'h97a217c1 ;
			32'h00100450 : data_o = 32'hfe87c803 ;
			32'h00100454 : data_o = 32'h17c177f9 ;
			32'h00100458 : data_o = 32'hc88397a2 ;
			32'h0010045c : data_o = 32'h4785fe87 ;
			32'h00100460 : data_o = 32'h879ac03e ;
			32'h00100464 : data_o = 32'h2e23339d ;
			32'h00100468 : data_o = 32'h2503fca4 ;
			32'h0010046c : data_o = 32'h35bdfdc4 ;
			32'h00100470 : data_o = 32'h853e4781 ;
			32'h00100474 : data_o = 32'h91166289 ;
			32'h00100478 : data_o = 32'h546250f2 ;
			32'h0010047c : data_o = 32'h80826121 ;
			32'h00100480 : data_o = 32'hd6067179 ;
			32'h00100484 : data_o = 32'h1800d422 ;
			32'h00100488 : data_o = 32'h0fa387aa ;
			32'h0010048c : data_o = 32'h4783fcf4 ;
			32'h00100490 : data_o = 32'h05a3fdf4 ;
			32'h00100494 : data_o = 32'h2623fef4 ;
			32'h00100498 : data_o = 32'ha835fe04 ;
			32'h0010049c : data_o = 32'hfeb44703 ;
			32'h001004a0 : data_o = 32'h77b347a9 ;
			32'h001004a4 : data_o = 32'hf79302f7 ;
			32'h001004a8 : data_o = 32'h87930ff7 ;
			32'h001004ac : data_o = 32'hf7130307 ;
			32'h001004b0 : data_o = 32'h27830ff7 ;
			32'h001004b4 : data_o = 32'h17c1fec4 ;
			32'h001004b8 : data_o = 32'h8a2397a2 ;
			32'h001004bc : data_o = 32'h4703fee7 ;
			32'h001004c0 : data_o = 32'h47a9feb4 ;
			32'h001004c4 : data_o = 32'h02f757b3 ;
			32'h001004c8 : data_o = 32'hfef405a3 ;
			32'h001004cc : data_o = 32'hfec42783 ;
			32'h001004d0 : data_o = 32'h26230785 ;
			32'h001004d4 : data_o = 32'h2703fef4 ;
			32'h001004d8 : data_o = 32'h478dfec4 ;
			32'h001004dc : data_o = 32'hfce7d0e3 ;
			32'h001004e0 : data_o = 32'h2623478d ;
			32'h001004e4 : data_o = 32'ha831fef4 ;
			32'h001004e8 : data_o = 32'hfec42783 ;
			32'h001004ec : data_o = 32'h97a217c1 ;
			32'h001004f0 : data_o = 32'hff47c783 ;
			32'h001004f4 : data_o = 32'h2aa9853e ;
			32'h001004f8 : data_o = 32'hfec42783 ;
			32'h001004fc : data_o = 32'h262317fd ;
			32'h00100500 : data_o = 32'h2783fef4 ;
			32'h00100504 : data_o = 32'hd1e3fec4 ;
			32'h00100508 : data_o = 32'h0001fe07 ;
			32'h0010050c : data_o = 32'h50b20001 ;
			32'h00100510 : data_o = 32'h61455422 ;
			32'h00100514 : data_o = 32'h715d8082 ;
			32'h00100518 : data_o = 32'hc4a2c686 ;
			32'h0010051c : data_o = 32'h0880c2a6 ;
			32'h00100520 : data_o = 32'hfaa42e23 ;
			32'h00100524 : data_o = 32'hfe0407a3 ;
			32'h00100528 : data_o = 32'h4783a881 ;
			32'h0010052c : data_o = 32'h8385fef4 ;
			32'h00100530 : data_o = 32'h0ff7f693 ;
			32'h00100534 : data_o = 32'hfbc42783 ;
			32'h00100538 : data_o = 32'h0ff7f593 ;
			32'h0010053c : data_o = 32'hfef44783 ;
			32'h00100540 : data_o = 32'h00178713 ;
			32'h00100544 : data_o = 32'h41f75793 ;
			32'h00100548 : data_o = 32'h973e83fd ;
			32'h0010054c : data_o = 32'h07b38b05 ;
			32'h00100550 : data_o = 32'hf79340f7 ;
			32'h00100554 : data_o = 32'h44830ff7 ;
			32'h00100558 : data_o = 32'h863efef4 ;
			32'h0010055c : data_o = 32'h33358536 ;
			32'h00100560 : data_o = 32'h9793872a ;
			32'h00100564 : data_o = 32'h17c10024 ;
			32'h00100568 : data_o = 32'hac2397a2 ;
			32'h0010056c : data_o = 32'h4783fce7 ;
			32'h00100570 : data_o = 32'h0785fef4 ;
			32'h00100574 : data_o = 32'hfef407a3 ;
			32'h00100578 : data_o = 32'hfef44703 ;
			32'h0010057c : data_o = 32'hf6e3479d ;
			32'h00100580 : data_o = 32'h07a3fae7 ;
			32'h00100584 : data_o = 32'ha095fe04 ;
			32'h00100588 : data_o = 32'hfef44783 ;
			32'h0010058c : data_o = 32'hf7938b85 ;
			32'h00100590 : data_o = 32'he7990ff7 ;
			32'h00100594 : data_o = 32'h02000513 ;
			32'h00100598 : data_o = 32'h05132865 ;
			32'h0010059c : data_o = 32'h284d07c0 ;
			32'h001005a0 : data_o = 32'h2423478d ;
			32'h001005a4 : data_o = 32'ha80dfef4 ;
			32'h001005a8 : data_o = 32'hfef44783 ;
			32'h001005ac : data_o = 32'h17c1078a ;
			32'h001005b0 : data_o = 32'ha70397a2 ;
			32'h001005b4 : data_o = 32'h2783fd87 ;
			32'h001005b8 : data_o = 32'h078efe84 ;
			32'h001005bc : data_o = 32'h00f757b3 ;
			32'h001005c0 : data_o = 32'h0ff7f793 ;
			32'h001005c4 : data_o = 32'h3d6d853e ;
			32'h001005c8 : data_o = 32'h07c00513 ;
			32'h001005cc : data_o = 32'h27832051 ;
			32'h001005d0 : data_o = 32'h17fdfe84 ;
			32'h001005d4 : data_o = 32'hfef42423 ;
			32'h001005d8 : data_o = 32'hfe842783 ;
			32'h001005dc : data_o = 32'hfc07d6e3 ;
			32'h001005e0 : data_o = 32'hfef44783 ;
			32'h001005e4 : data_o = 32'h07a30785 ;
			32'h001005e8 : data_o = 32'h4703fef4 ;
			32'h001005ec : data_o = 32'h479dfef4 ;
			32'h001005f0 : data_o = 32'hf8e7fce3 ;
			32'h001005f4 : data_o = 32'h02000513 ;
			32'h001005f8 : data_o = 32'h452928a1 ;
			32'h001005fc : data_o = 32'h00012891 ;
			32'h00100600 : data_o = 32'h442640b6 ;
			32'h00100604 : data_o = 32'h61614496 ;
			32'h00100608 : data_o = 32'h11018082 ;
			32'h0010060c : data_o = 32'hcc22ce06 ;
			32'h00100610 : data_o = 32'h26231000 ;
			32'h00100614 : data_o = 32'ha00dfe04 ;
			32'h00100618 : data_o = 32'hfec42783 ;
			32'h0010061c : data_o = 32'h03f7f793 ;
			32'h00100620 : data_o = 32'h4529e399 ;
			32'h00100624 : data_o = 32'h27832035 ;
			32'h00100628 : data_o = 32'h853efec4 ;
			32'h0010062c : data_o = 32'h278335ed ;
			32'h00100630 : data_o = 32'h0785fec4 ;
			32'h00100634 : data_o = 32'hfef42623 ;
			32'h00100638 : data_o = 32'hfec42703 ;
			32'h0010063c : data_o = 32'h1ff00793 ;
			32'h00100640 : data_o = 32'hfce7dce3 ;
			32'h00100644 : data_o = 32'h00010001 ;
			32'h00100648 : data_o = 32'h446240f2 ;
			32'h0010064c : data_o = 32'h80826105 ;
			32'h00100650 : data_o = 32'hce221101 ;
			32'h00100654 : data_o = 32'h87aa1000 ;
			32'h00100658 : data_o = 32'hfef407a3 ;
			32'h0010065c : data_o = 32'h000207b7 ;
			32'h00100660 : data_o = 32'hfef44703 ;
			32'h00100664 : data_o = 32'h4783c398 ;
			32'h00100668 : data_o = 32'h853efef4 ;
			32'h0010066c : data_o = 32'h61054472 ;
			32'h00100670 : data_o = 32'h11418082 ;
			32'h00100674 : data_o = 32'hc422c606 ;
			32'h00100678 : data_o = 32'h15370800 ;
			32'h0010067c : data_o = 32'h24c58000 ;
			32'h00100680 : data_o = 32'h853e87aa ;
			32'h00100684 : data_o = 32'h442240b2 ;
			32'h00100688 : data_o = 32'h80820141 ;
			32'h0010068c : data_o = 32'hce061101 ;
			32'h00100690 : data_o = 32'h1000cc22 ;
			32'h00100694 : data_o = 32'hfea42623 ;
			32'h00100698 : data_o = 32'h2783a819 ;
			32'h0010069c : data_o = 32'h8713fec4 ;
			32'h001006a0 : data_o = 32'h26230017 ;
			32'h001006a4 : data_o = 32'hc783fee4 ;
			32'h001006a8 : data_o = 32'h853e0007 ;
			32'h001006ac : data_o = 32'h27833755 ;
			32'h001006b0 : data_o = 32'hc783fec4 ;
			32'h001006b4 : data_o = 32'hf3f50007 ;
			32'h001006b8 : data_o = 32'h853e4781 ;
			32'h001006bc : data_o = 32'h446240f2 ;
			32'h001006c0 : data_o = 32'h80826105 ;
			32'h001006c4 : data_o = 32'hd6067179 ;
			32'h001006c8 : data_o = 32'h1800d422 ;
			32'h001006cc : data_o = 32'hfca42e23 ;
			32'h001006d0 : data_o = 32'hfe042623 ;
			32'h001006d4 : data_o = 32'h2783a891 ;
			32'h001006d8 : data_o = 32'h83f1fdc4 ;
			32'h001006dc : data_o = 32'hfef42423 ;
			32'h001006e0 : data_o = 32'hfe842703 ;
			32'h001006e4 : data_o = 32'hcd6347a5 ;
			32'h001006e8 : data_o = 32'h278300e7 ;
			32'h001006ec : data_o = 32'hf793fe84 ;
			32'h001006f0 : data_o = 32'h87930ff7 ;
			32'h001006f4 : data_o = 32'hf7930307 ;
			32'h001006f8 : data_o = 32'h853e0ff7 ;
			32'h001006fc : data_o = 32'ha8193f91 ;
			32'h00100700 : data_o = 32'hfe842783 ;
			32'h00100704 : data_o = 32'h0ff7f793 ;
			32'h00100708 : data_o = 32'h03778793 ;
			32'h0010070c : data_o = 32'h0ff7f793 ;
			32'h00100710 : data_o = 32'h3f3d853e ;
			32'h00100714 : data_o = 32'hfdc42783 ;
			32'h00100718 : data_o = 32'h2e230792 ;
			32'h0010071c : data_o = 32'h2783fcf4 ;
			32'h00100720 : data_o = 32'h0785fec4 ;
			32'h00100724 : data_o = 32'hfef42623 ;
			32'h00100728 : data_o = 32'hfec42703 ;
			32'h0010072c : data_o = 32'hd4e3479d ;
			32'h00100730 : data_o = 32'h0001fae7 ;
			32'h00100734 : data_o = 32'h50b20001 ;
			32'h00100738 : data_o = 32'h61455422 ;
			32'h0010073c : data_o = 32'h11418082 ;
			32'h00100740 : data_o = 32'h0800c622 ;
			32'h00100744 : data_o = 32'h000207b7 ;
			32'h00100748 : data_o = 32'h470507a1 ;
			32'h0010074c : data_o = 32'h0001c398 ;
			32'h00100750 : data_o = 32'h01414432 ;
			32'h00100754 : data_o = 32'h11018082 ;
			32'h00100758 : data_o = 32'h1000ce22 ;
			32'h0010075c : data_o = 32'h341027f3 ;
			32'h00100760 : data_o = 32'hfef42623 ;
			32'h00100764 : data_o = 32'hfec42783 ;
			32'h00100768 : data_o = 32'h4472853e ;
			32'h0010076c : data_o = 32'h80826105 ;
			32'h00100770 : data_o = 32'hce221101 ;
			32'h00100774 : data_o = 32'h27f31000 ;
			32'h00100778 : data_o = 32'h26233420 ;
			32'h0010077c : data_o = 32'h2783fef4 ;
			32'h00100780 : data_o = 32'h853efec4 ;
			32'h00100784 : data_o = 32'h61054472 ;
			32'h00100788 : data_o = 32'h11018082 ;
			32'h0010078c : data_o = 32'h1000ce22 ;
			32'h00100790 : data_o = 32'h343027f3 ;
			32'h00100794 : data_o = 32'hfef42623 ;
			32'h00100798 : data_o = 32'hfec42783 ;
			32'h0010079c : data_o = 32'h4472853e ;
			32'h001007a0 : data_o = 32'h80826105 ;
			32'h001007a4 : data_o = 32'hce221101 ;
			32'h001007a8 : data_o = 32'h27f31000 ;
			32'h001007ac : data_o = 32'h2623b000 ;
			32'h001007b0 : data_o = 32'h2783fef4 ;
			32'h001007b4 : data_o = 32'h853efec4 ;
			32'h001007b8 : data_o = 32'h61054472 ;
			32'h001007bc : data_o = 32'h11418082 ;
			32'h001007c0 : data_o = 32'h0800c622 ;
			32'h001007c4 : data_o = 32'hb0001073 ;
			32'h001007c8 : data_o = 32'h44320001 ;
			32'h001007cc : data_o = 32'h80820141 ;
			32'h001007d0 : data_o = 32'hd6227179 ;
			32'h001007d4 : data_o = 32'h2e231800 ;
			32'h001007d8 : data_o = 32'h2c23fca4 ;
			32'h001007dc : data_o = 32'h2703fcb4 ;
			32'h001007e0 : data_o = 32'h47fdfdc4 ;
			32'h001007e4 : data_o = 32'h00e7f463 ;
			32'h001007e8 : data_o = 32'ha8794785 ;
			32'h001007ec : data_o = 32'h00100797 ;
			32'h001007f0 : data_o = 32'h81478793 ;
			32'h001007f4 : data_o = 32'h27834398 ;
			32'h001007f8 : data_o = 32'h078afdc4 ;
			32'h001007fc : data_o = 32'h262397ba ;
			32'h00100800 : data_o = 32'h2703fef4 ;
			32'h00100804 : data_o = 32'h2783fd84 ;
			32'h00100808 : data_o = 32'h07b3fec4 ;
			32'h0010080c : data_o = 32'h242340f7 ;
			32'h00100810 : data_o = 32'h2703fef4 ;
			32'h00100814 : data_o = 32'h07b7fe84 ;
			32'h00100818 : data_o = 32'h58630008 ;
			32'h0010081c : data_o = 32'h270300f7 ;
			32'h00100820 : data_o = 32'h07b7fe84 ;
			32'h00100824 : data_o = 32'h5463fff8 ;
			32'h00100828 : data_o = 32'h478900f7 ;
			32'h0010082c : data_o = 32'h2783a8b1 ;
			32'h00100830 : data_o = 32'h2223fe84 ;
			32'h00100834 : data_o = 32'h2783fef4 ;
			32'h00100838 : data_o = 32'h9713fe44 ;
			32'h0010083c : data_o = 32'h07b70147 ;
			32'h00100840 : data_o = 32'h8f7d7fe0 ;
			32'h00100844 : data_o = 32'hfe442783 ;
			32'h00100848 : data_o = 32'h00979693 ;
			32'h0010084c : data_o = 32'h001007b7 ;
			32'h00100850 : data_o = 32'h8f5d8ff5 ;
			32'h00100854 : data_o = 32'hfe442683 ;
			32'h00100858 : data_o = 32'h000ff7b7 ;
			32'h0010085c : data_o = 32'h8f5d8ff5 ;
			32'h00100860 : data_o = 32'hfe442783 ;
			32'h00100864 : data_o = 32'h00b79693 ;
			32'h00100868 : data_o = 32'h800007b7 ;
			32'h0010086c : data_o = 32'h8fd98ff5 ;
			32'h00100870 : data_o = 32'h06f7e793 ;
			32'h00100874 : data_o = 32'hfef42023 ;
			32'h00100878 : data_o = 32'hfec42783 ;
			32'h0010087c : data_o = 32'hfe042703 ;
			32'h00100880 : data_o = 32'h100fc398 ;
			32'h00100884 : data_o = 32'h47810000 ;
			32'h00100888 : data_o = 32'h5432853e ;
			32'h0010088c : data_o = 32'h80826145 ;
			32'h00100890 : data_o = 32'hce221101 ;
			32'h00100894 : data_o = 32'h26231000 ;
			32'h00100898 : data_o = 32'h2783fea4 ;
			32'h0010089c : data_o = 32'ha073fec4 ;
			32'h001008a0 : data_o = 32'h00013047 ;
			32'h001008a4 : data_o = 32'h61054472 ;
			32'h001008a8 : data_o = 32'h11018082 ;
			32'h001008ac : data_o = 32'h1000ce22 ;
			32'h001008b0 : data_o = 32'hfea42623 ;
			32'h001008b4 : data_o = 32'hfec42783 ;
			32'h001008b8 : data_o = 32'h3047b073 ;
			32'h001008bc : data_o = 32'h44720001 ;
			32'h001008c0 : data_o = 32'h80826105 ;
			32'h001008c4 : data_o = 32'hce221101 ;
			32'h001008c8 : data_o = 32'h26231000 ;
			32'h001008cc : data_o = 32'h2783fea4 ;
			32'h001008d0 : data_o = 32'hc789fec4 ;
			32'h001008d4 : data_o = 32'ha07347a1 ;
			32'h001008d8 : data_o = 32'ha0213007 ;
			32'h001008dc : data_o = 32'hb07347a1 ;
			32'h001008e0 : data_o = 32'h00013007 ;
			32'h001008e4 : data_o = 32'h61054472 ;
			32'h001008e8 : data_o = 32'h11418082 ;
			32'h001008ec : data_o = 32'hc422c606 ;
			32'h001008f0 : data_o = 32'h25170800 ;
			32'h001008f4 : data_o = 32'h05130000 ;
			32'h001008f8 : data_o = 32'h3b497965 ;
			32'h001008fc : data_o = 32'h00002517 ;
			32'h00100900 : data_o = 32'h79c50513 ;
			32'h00100904 : data_o = 32'h25173361 ;
			32'h00100908 : data_o = 32'h05130000 ;
			32'h0010090c : data_o = 32'h3bbd7a25 ;
			32'h00100910 : data_o = 32'h87aa3599 ;
			32'h00100914 : data_o = 32'h337d853e ;
			32'h00100918 : data_o = 32'h00002517 ;
			32'h0010091c : data_o = 32'h79c50513 ;
			32'h00100920 : data_o = 32'h35b933b5 ;
			32'h00100924 : data_o = 32'h853e87aa ;
			32'h00100928 : data_o = 32'h25173b71 ;
			32'h0010092c : data_o = 32'h05130000 ;
			32'h00100930 : data_o = 32'h3ba97965 ;
			32'h00100934 : data_o = 32'h87aa3d99 ;
			32'h00100938 : data_o = 32'h3369853e ;
			32'h0010093c : data_o = 32'h3b094529 ;
			32'h00100940 : data_o = 32'hbffd0001 ;
			32'h00100944 : data_o = 32'hc6061141 ;
			32'h00100948 : data_o = 32'h0800c422 ;
			32'h0010094c : data_o = 32'h37896541 ;
			32'h00100950 : data_o = 32'h3f8d4505 ;
			32'h00100954 : data_o = 32'h40b20001 ;
			32'h00100958 : data_o = 32'h01414422 ;
			32'h0010095c : data_o = 32'h71798082 ;
			32'h00100960 : data_o = 32'h1800d622 ;
			32'h00100964 : data_o = 32'hfca42e23 ;
			32'h00100968 : data_o = 32'h262357fd ;
			32'h0010096c : data_o = 32'h2783fef4 ;
			32'h00100970 : data_o = 32'h07a1fdc4 ;
			32'h00100974 : data_o = 32'h8b85439c ;
			32'h00100978 : data_o = 32'h2783e791 ;
			32'h0010097c : data_o = 32'h439cfdc4 ;
			32'h00100980 : data_o = 32'hfef42623 ;
			32'h00100984 : data_o = 32'hfec42783 ;
			32'h00100988 : data_o = 32'h5432853e ;
			32'h0010098c : data_o = 32'h80826145 ;
			32'h00100990 : data_o = 32'hce221101 ;
			32'h00100994 : data_o = 32'h26231000 ;
			32'h00100998 : data_o = 32'h87aefea4 ;
			32'h0010099c : data_o = 32'hfef405a3 ;
			32'h001009a0 : data_o = 32'h27830001 ;
			32'h001009a4 : data_o = 32'h07a1fec4 ;
			32'h001009a8 : data_o = 32'h8b89439c ;
			32'h001009ac : data_o = 32'h2783fbfd ;
			32'h001009b0 : data_o = 32'h0791fec4 ;
			32'h001009b4 : data_o = 32'hfeb44703 ;
			32'h001009b8 : data_o = 32'h0001c398 ;
			32'h001009bc : data_o = 32'h61054472 ;
			32'h001009c0 : data_o = 32'h11018082 ;
			32'h001009c4 : data_o = 32'h1000ce22 ;
			32'h001009c8 : data_o = 32'hfea42423 ;
			32'h001009cc : data_o = 32'hfeb42623 ;
			32'h001009d0 : data_o = 32'h080026b7 ;
			32'h001009d4 : data_o = 32'h567d06a1 ;
			32'h001009d8 : data_o = 32'h2683c290 ;
			32'h001009dc : data_o = 32'hd713fec4 ;
			32'h001009e0 : data_o = 32'h47810006 ;
			32'h001009e4 : data_o = 32'h080026b7 ;
			32'h001009e8 : data_o = 32'h87ba06b1 ;
			32'h001009ec : data_o = 32'h27b7c29c ;
			32'h001009f0 : data_o = 32'h07a10800 ;
			32'h001009f4 : data_o = 32'hfe842703 ;
			32'h001009f8 : data_o = 32'h0001c398 ;
			32'h001009fc : data_o = 32'h61054472 ;
			32'h00100a00 : data_o = 32'h71798082 ;
			32'h00100a04 : data_o = 32'hd422d606 ;
			32'h00100a08 : data_o = 32'h2c231800 ;
			32'h00100a0c : data_o = 32'h2e23fca4 ;
			32'h00100a10 : data_o = 32'h20fdfcb4 ;
			32'h00100a14 : data_o = 32'hfea42423 ;
			32'h00100a18 : data_o = 32'hfeb42623 ;
			32'h00100a1c : data_o = 32'hfe842603 ;
			32'h00100a20 : data_o = 32'hfec42683 ;
			32'h00100a24 : data_o = 32'hfd842503 ;
			32'h00100a28 : data_o = 32'hfdc42583 ;
			32'h00100a2c : data_o = 32'h00a60733 ;
			32'h00100a30 : data_o = 32'h3833883a ;
			32'h00100a34 : data_o = 32'h87b300c8 ;
			32'h00100a38 : data_o = 32'h06b300b6 ;
			32'h00100a3c : data_o = 32'h87b600f8 ;
			32'h00100a40 : data_o = 32'hfee42423 ;
			32'h00100a44 : data_o = 32'hfef42623 ;
			32'h00100a48 : data_o = 32'hfe842503 ;
			32'h00100a4c : data_o = 32'hfec42583 ;
			32'h00100a50 : data_o = 32'h00013f8d ;
			32'h00100a54 : data_o = 32'h542250b2 ;
			32'h00100a58 : data_o = 32'h80826145 ;
			32'h00100a5c : data_o = 32'hc686715d ;
			32'h00100a60 : data_o = 32'hc29ac496 ;
			32'h00100a64 : data_o = 32'hde22c09e ;
			32'h00100a68 : data_o = 32'hda2edc2a ;
			32'h00100a6c : data_o = 32'hd636d832 ;
			32'h00100a70 : data_o = 32'hd23ed43a ;
			32'h00100a74 : data_o = 32'hce46d042 ;
			32'h00100a78 : data_o = 32'hca76cc72 ;
			32'h00100a7c : data_o = 32'hc67ec87a ;
			32'h00100a80 : data_o = 32'hf7970880 ;
			32'h00100a84 : data_o = 32'h8793000f ;
			32'h00100a88 : data_o = 32'h43985a67 ;
			32'h00100a8c : data_o = 32'h853a43dc ;
			32'h00100a90 : data_o = 32'h3f8585be ;
			32'h00100a94 : data_o = 32'h000ff797 ;
			32'h00100a98 : data_o = 32'h58c78793 ;
			32'h00100a9c : data_o = 32'h43dc4398 ;
			32'h00100aa0 : data_o = 32'h45814505 ;
			32'h00100aa4 : data_o = 32'h00a70633 ;
			32'h00100aa8 : data_o = 32'h38338832 ;
			32'h00100aac : data_o = 32'h86b300e8 ;
			32'h00100ab0 : data_o = 32'h07b300b7 ;
			32'h00100ab4 : data_o = 32'h86be00d8 ;
			32'h00100ab8 : data_o = 32'h87b68732 ;
			32'h00100abc : data_o = 32'h000ff697 ;
			32'h00100ac0 : data_o = 32'h56468693 ;
			32'h00100ac4 : data_o = 32'hc2dcc298 ;
			32'h00100ac8 : data_o = 32'h40b60001 ;
			32'h00100acc : data_o = 32'h431642a6 ;
			32'h00100ad0 : data_o = 32'h54724386 ;
			32'h00100ad4 : data_o = 32'h55d25562 ;
			32'h00100ad8 : data_o = 32'h56b25642 ;
			32'h00100adc : data_o = 32'h57925722 ;
			32'h00100ae0 : data_o = 32'h48f25802 ;
			32'h00100ae4 : data_o = 32'h4ed24e62 ;
			32'h00100ae8 : data_o = 32'h4fb24f42 ;
			32'h00100aec : data_o = 32'h00736161 ;
			32'h00100af0 : data_o = 32'h11413020 ;
			32'h00100af4 : data_o = 32'h0800c622 ;
			32'h00100af8 : data_o = 32'h44320001 ;
			32'h00100afc : data_o = 32'h80820141 ;
			32'h00100b00 : data_o = 32'hce221101 ;
			32'h00100b04 : data_o = 32'h28371000 ;
			32'h00100b08 : data_o = 32'h08110800 ;
			32'h00100b0c : data_o = 32'h00082803 ;
			32'h00100b10 : data_o = 32'hff042623 ;
			32'h00100b14 : data_o = 32'h08002837 ;
			32'h00100b18 : data_o = 32'h00082803 ;
			32'h00100b1c : data_o = 32'hff042423 ;
			32'h00100b20 : data_o = 32'h08002837 ;
			32'h00100b24 : data_o = 32'h28030811 ;
			32'h00100b28 : data_o = 32'h28830008 ;
			32'h00100b2c : data_o = 32'h9ce3fec4 ;
			32'h00100b30 : data_o = 32'h2803fd08 ;
			32'h00100b34 : data_o = 32'h8542fec4 ;
			32'h00100b38 : data_o = 32'h17934581 ;
			32'h00100b3c : data_o = 32'h47010005 ;
			32'h00100b40 : data_o = 32'hfe842583 ;
			32'h00100b44 : data_o = 32'h4681862e ;
			32'h00100b48 : data_o = 32'h00c765b3 ;
			32'h00100b4c : data_o = 32'hfeb42023 ;
			32'h00100b50 : data_o = 32'h22238fd5 ;
			32'h00100b54 : data_o = 32'h2703fef4 ;
			32'h00100b58 : data_o = 32'h2783fe04 ;
			32'h00100b5c : data_o = 32'h853afe44 ;
			32'h00100b60 : data_o = 32'h447285be ;
			32'h00100b64 : data_o = 32'h80826105 ;
			32'h00100b68 : data_o = 32'hc6221141 ;
			32'h00100b6c : data_o = 32'hf7970800 ;
			32'h00100b70 : data_o = 32'h8793000f ;
			32'h00100b74 : data_o = 32'h43984b27 ;
			32'h00100b78 : data_o = 32'h853a43dc ;
			32'h00100b7c : data_o = 32'h443285be ;
			32'h00100b80 : data_o = 32'h80820141 ;
			32'h00100b84 : data_o = 32'hce061101 ;
			32'h00100b88 : data_o = 32'h1000cc22 ;
			32'h00100b8c : data_o = 32'hfea42423 ;
			32'h00100b90 : data_o = 32'hfeb42623 ;
			32'h00100b94 : data_o = 32'h000ff797 ;
			32'h00100b98 : data_o = 32'h48c78793 ;
			32'h00100b9c : data_o = 32'h47014681 ;
			32'h00100ba0 : data_o = 32'hc3d8c394 ;
			32'h00100ba4 : data_o = 32'h000ff697 ;
			32'h00100ba8 : data_o = 32'h48468693 ;
			32'h00100bac : data_o = 32'hfe842703 ;
			32'h00100bb0 : data_o = 32'hfec42783 ;
			32'h00100bb4 : data_o = 32'hc2dcc298 ;
			32'h00100bb8 : data_o = 32'hfe842503 ;
			32'h00100bbc : data_o = 32'hfec42583 ;
			32'h00100bc0 : data_o = 32'h05133589 ;
			32'h00100bc4 : data_o = 32'h31e90800 ;
			32'h00100bc8 : data_o = 32'h39ed4505 ;
			32'h00100bcc : data_o = 32'h40f20001 ;
			32'h00100bd0 : data_o = 32'h61054462 ;
			32'h00100bd4 : data_o = 32'h11418082 ;
			32'h00100bd8 : data_o = 32'h0800c622 ;
			32'h00100bdc : data_o = 32'h08000793 ;
			32'h00100be0 : data_o = 32'h3047b073 ;
			32'h00100be4 : data_o = 32'h44320001 ;
			32'h00100be8 : data_o = 32'h80820141 ;
			32'h00100bec : data_o = 32'hce221101 ;
			32'h00100bf0 : data_o = 32'h26231000 ;
			32'h00100bf4 : data_o = 32'h2423fea4 ;
			32'h00100bf8 : data_o = 32'h2783feb4 ;
			32'h00100bfc : data_o = 32'h2703fec4 ;
			32'h00100c00 : data_o = 32'hc398fe84 ;
			32'h00100c04 : data_o = 32'h44720001 ;
			32'h00100c08 : data_o = 32'h80826105 ;
			32'h00100c0c : data_o = 32'hce221101 ;
			32'h00100c10 : data_o = 32'h26231000 ;
			32'h00100c14 : data_o = 32'h2783fea4 ;
			32'h00100c18 : data_o = 32'h439cfec4 ;
			32'h00100c1c : data_o = 32'h4472853e ;
			32'h00100c20 : data_o = 32'h80826105 ;
			32'h00100c24 : data_o = 32'hd6067179 ;
			32'h00100c28 : data_o = 32'h1800d422 ;
			32'h00100c2c : data_o = 32'hfca42e23 ;
			32'h00100c30 : data_o = 32'hfcb42c23 ;
			32'h00100c34 : data_o = 32'hfcc42a23 ;
			32'h00100c38 : data_o = 32'hfdc42503 ;
			32'h00100c3c : data_o = 32'h26233fc1 ;
			32'h00100c40 : data_o = 32'h2783fea4 ;
			32'h00100c44 : data_o = 32'h4705fd84 ;
			32'h00100c48 : data_o = 32'h00f717b3 ;
			32'h00100c4c : data_o = 32'hfff7c793 ;
			32'h00100c50 : data_o = 32'h2783873e ;
			32'h00100c54 : data_o = 32'h8ff9fec4 ;
			32'h00100c58 : data_o = 32'hfef42623 ;
			32'h00100c5c : data_o = 32'hfd842783 ;
			32'h00100c60 : data_o = 32'hfd442703 ;
			32'h00100c64 : data_o = 32'h00f717b3 ;
			32'h00100c68 : data_o = 32'hfec42703 ;
			32'h00100c6c : data_o = 32'h26238fd9 ;
			32'h00100c70 : data_o = 32'h2583fef4 ;
			32'h00100c74 : data_o = 32'h2503fec4 ;
			32'h00100c78 : data_o = 32'h3f8dfdc4 ;
			32'h00100c7c : data_o = 32'h50b20001 ;
			32'h00100c80 : data_o = 32'h61455422 ;
			32'h00100c84 : data_o = 32'h71798082 ;
			32'h00100c88 : data_o = 32'hd422d606 ;
			32'h00100c8c : data_o = 32'h2e231800 ;
			32'h00100c90 : data_o = 32'h2c23fca4 ;
			32'h00100c94 : data_o = 32'h2503fcb4 ;
			32'h00100c98 : data_o = 32'h3f8dfdc4 ;
			32'h00100c9c : data_o = 32'hfea42623 ;
			32'h00100ca0 : data_o = 32'hfd842783 ;
			32'h00100ca4 : data_o = 32'hfec42703 ;
			32'h00100ca8 : data_o = 32'h00f757b3 ;
			32'h00100cac : data_o = 32'h853e8b85 ;
			32'h00100cb0 : data_o = 32'h542250b2 ;
			32'h00100cb4 : data_o = 32'h80826145 ;
			32'h00100cb8 : data_o = 32'hce221101 ;
			32'h00100cbc : data_o = 32'h26231000 ;
			32'h00100cc0 : data_o = 32'h07b7fea4 ;
			32'h00100cc4 : data_o = 32'h07c17000 ;
			32'h00100cc8 : data_o = 32'hfec42703 ;
			32'h00100ccc : data_o = 32'h0001c398 ;
			32'h00100cd0 : data_o = 32'h61054472 ;
			32'h00100cd4 : data_o = 32'h71798082 ;
			32'h00100cd8 : data_o = 32'h1800d622 ;
			32'h00100cdc : data_o = 32'h873687aa ;
			32'h00100ce0 : data_o = 32'hfcf40fa3 ;
			32'h00100ce4 : data_o = 32'h0f2387ae ;
			32'h00100ce8 : data_o = 32'h87b2fcf4 ;
			32'h00100cec : data_o = 32'hfcf40ea3 ;
			32'h00100cf0 : data_o = 32'h0e2387ba ;
			32'h00100cf4 : data_o = 32'h4703fcf4 ;
			32'h00100cf8 : data_o = 32'h4783fdf4 ;
			32'h00100cfc : data_o = 32'h07a2fde4 ;
			32'h00100d00 : data_o = 32'h47838f5d ;
			32'h00100d04 : data_o = 32'h07c2fdd4 ;
			32'h00100d08 : data_o = 32'h47838f5d ;
			32'h00100d0c : data_o = 32'h07e2fdc4 ;
			32'h00100d10 : data_o = 32'h26238fd9 ;
			32'h00100d14 : data_o = 32'h07b7fef4 ;
			32'h00100d18 : data_o = 32'h87937000 ;
			32'h00100d1c : data_o = 32'h27030347 ;
			32'h00100d20 : data_o = 32'hc398fec4 ;
			32'h00100d24 : data_o = 32'h54320001 ;
			32'h00100d28 : data_o = 32'h80826145 ;
			32'h00100d2c : data_o = 32'hd6227179 ;
			32'h00100d30 : data_o = 32'h87aa1800 ;
			32'h00100d34 : data_o = 32'h0fa38736 ;
			32'h00100d38 : data_o = 32'h87aefcf4 ;
			32'h00100d3c : data_o = 32'hfcf40f23 ;
			32'h00100d40 : data_o = 32'h0ea387b2 ;
			32'h00100d44 : data_o = 32'h87bafcf4 ;
			32'h00100d48 : data_o = 32'hfcf40e23 ;
			32'h00100d4c : data_o = 32'hfdf44703 ;
			32'h00100d50 : data_o = 32'hfde44783 ;
			32'h00100d54 : data_o = 32'h8f5d07a2 ;
			32'h00100d58 : data_o = 32'hfdd44783 ;
			32'h00100d5c : data_o = 32'h8f5d07c2 ;
			32'h00100d60 : data_o = 32'hfdc44783 ;
			32'h00100d64 : data_o = 32'h8fd907e2 ;
			32'h00100d68 : data_o = 32'hfef42623 ;
			32'h00100d6c : data_o = 32'h700007b7 ;
			32'h00100d70 : data_o = 32'h03878793 ;
			32'h00100d74 : data_o = 32'hfec42703 ;
			32'h00100d78 : data_o = 32'h0001c398 ;
			32'h00100d7c : data_o = 32'h61455432 ;
			32'h00100d80 : data_o = 32'h11018082 ;
			32'h00100d84 : data_o = 32'h1000ce22 ;
			32'h00100d88 : data_o = 32'hfea42623 ;
			32'h00100d8c : data_o = 32'h700007b7 ;
			32'h00100d90 : data_o = 32'h02078793 ;
			32'h00100d94 : data_o = 32'hfec42703 ;
			32'h00100d98 : data_o = 32'h0001c398 ;
			32'h00100d9c : data_o = 32'h61054472 ;
			32'h00100da0 : data_o = 32'h11418082 ;
			32'h00100da4 : data_o = 32'h0800c622 ;
			32'h00100da8 : data_o = 32'h700007b7 ;
			32'h00100dac : data_o = 32'h02478793 ;
			32'h00100db0 : data_o = 32'hc3984705 ;
			32'h00100db4 : data_o = 32'h44320001 ;
			32'h00100db8 : data_o = 32'h80820141 ;
			32'h00100dbc : data_o = 32'hc6221141 ;
			32'h00100dc0 : data_o = 32'h07b70800 ;
			32'h00100dc4 : data_o = 32'h87937000 ;
			32'h00100dc8 : data_o = 32'h439c0287 ;
			32'h00100dcc : data_o = 32'h4432853e ;
			32'h00100dd0 : data_o = 32'h80820141 ;
			32'h00100dd4 : data_o = 32'hc6221141 ;
			32'h00100dd8 : data_o = 32'h07b70800 ;
			32'h00100ddc : data_o = 32'h87937000 ;
			32'h00100de0 : data_o = 32'h439c02c7 ;
			32'h00100de4 : data_o = 32'h4432853e ;
			32'h00100de8 : data_o = 32'h80820141 ;
			32'h00100dec : data_o = 32'hc6221141 ;
			32'h00100df0 : data_o = 32'h07b70800 ;
			32'h00100df4 : data_o = 32'h87937000 ;
			32'h00100df8 : data_o = 32'h439c0307 ;
			32'h00100dfc : data_o = 32'h4432853e ;
			32'h00100e00 : data_o = 32'h80820141 ;
			32'h00100e04 : data_o = 32'hce221101 ;
			32'h00100e08 : data_o = 32'h26231000 ;
			32'h00100e0c : data_o = 32'h2703fea4 ;
			32'h00100e10 : data_o = 32'h07b7fec4 ;
			32'h00100e14 : data_o = 32'h87937000 ;
			32'h00100e18 : data_o = 32'h97ba1007 ;
			32'h00100e1c : data_o = 32'h853e439c ;
			32'h00100e20 : data_o = 32'h61054472 ;
			32'h00100e24 : data_o = 32'h11018082 ;
			32'h00100e28 : data_o = 32'h1000ce22 ;
			32'h00100e2c : data_o = 32'hfea42623 ;
			32'h00100e30 : data_o = 32'h700007b7 ;
			32'h00100e34 : data_o = 32'h270307e1 ;
			32'h00100e38 : data_o = 32'hc398fec4 ;
			32'h00100e3c : data_o = 32'h44720001 ;
			32'h00100e40 : data_o = 32'h80826105 ;
			32'h00100e44 : data_o = 32'hce221101 ;
			32'h00100e48 : data_o = 32'h26231000 ;
			32'h00100e4c : data_o = 32'h07b7fea4 ;
			32'h00100e50 : data_o = 32'h87937000 ;
			32'h00100e54 : data_o = 32'h270303c7 ;
			32'h00100e58 : data_o = 32'hc398fec4 ;
			32'h00100e5c : data_o = 32'h44720001 ;
			32'h00100e60 : data_o = 32'h80826105 ;
			32'h00100e64 : data_o = 32'hce221101 ;
			32'h00100e68 : data_o = 32'h26231000 ;
			32'h00100e6c : data_o = 32'h87aefea4 ;
			32'h00100e70 : data_o = 32'h05a38736 ;
			32'h00100e74 : data_o = 32'h87b2fef4 ;
			32'h00100e78 : data_o = 32'hfef40523 ;
			32'h00100e7c : data_o = 32'h04a387ba ;
			32'h00100e80 : data_o = 32'h4783fef4 ;
			32'h00100e84 : data_o = 32'h078efeb4 ;
			32'h00100e88 : data_o = 32'h0187f713 ;
			32'h00100e8c : data_o = 32'hfea44783 ;
			32'h00100e90 : data_o = 32'h8f5d0796 ;
			32'h00100e94 : data_o = 32'hfe944783 ;
			32'h00100e98 : data_o = 32'h8b91078a ;
			32'h00100e9c : data_o = 32'h07b78f5d ;
			32'h00100ea0 : data_o = 32'h87937000 ;
			32'h00100ea4 : data_o = 32'h97ba1007 ;
			32'h00100ea8 : data_o = 32'h2783873e ;
			32'h00100eac : data_o = 32'hc793fec4 ;
			32'h00100eb0 : data_o = 32'hc31cfff7 ;
			32'h00100eb4 : data_o = 32'h44720001 ;
			32'h00100eb8 : data_o = 32'h80826105 ;
			32'h00100ebc : data_o = 32'ha2fff06f ;
			32'h00100ec0 : data_o = 32'h00000093 ;
			32'h00100ec4 : data_o = 32'h81868106 ;
			32'h00100ec8 : data_o = 32'h82868206 ;
			32'h00100ecc : data_o = 32'h83868306 ;
			32'h00100ed0 : data_o = 32'h84868406 ;
			32'h00100ed4 : data_o = 32'h85868506 ;
			32'h00100ed8 : data_o = 32'h86868606 ;
			32'h00100edc : data_o = 32'h87868706 ;
			32'h00100ee0 : data_o = 32'h88868806 ;
			32'h00100ee4 : data_o = 32'h89868906 ;
			32'h00100ee8 : data_o = 32'h8a868a06 ;
			32'h00100eec : data_o = 32'h8b868b06 ;
			32'h00100ef0 : data_o = 32'h8c868c06 ;
			32'h00100ef4 : data_o = 32'h8d868d06 ;
			32'h00100ef8 : data_o = 32'h8e868e06 ;
			32'h00100efc : data_o = 32'h8f868f06 ;
			32'h00100f00 : data_o = 32'h0011f117 ;
			32'h00100f04 : data_o = 32'h10010113 ;
			32'h00100f08 : data_o = 32'h000ffd17 ;
			32'h00100f0c : data_o = 32'h100d0d13 ;
			32'h00100f10 : data_o = 32'h000ffd97 ;
			32'h00100f14 : data_o = 32'h120d8d93 ;
			32'h00100f18 : data_o = 32'h01bd5763 ;
			32'h00100f1c : data_o = 32'h000d2023 ;
			32'h00100f20 : data_o = 32'hdde30d11 ;
			32'h00100f24 : data_o = 32'h4501ffad ;
			32'h00100f28 : data_o = 32'hf0ef4581 ;
			32'h00100f2c : data_o = 32'h02b7c46f ;
			32'h00100f30 : data_o = 32'h02a10002 ;
			32'h00100f34 : data_o = 32'ha0234305 ;
			32'h00100f38 : data_o = 32'h00730062 ;
			32'h00100f3c : data_o = 32'hbff51050 ;
			32'h00100f40 : data_o = 32'h00b547b3 ;
			32'h00100f44 : data_o = 32'h08b38b8d ;
			32'h00100f48 : data_o = 32'he7b100c5 ;
			32'h00100f4c : data_o = 32'hf463478d ;
			32'h00100f50 : data_o = 32'h779304c7 ;
			32'h00100f54 : data_o = 32'h872a0035 ;
			32'h00100f58 : data_o = 32'hf613ebb9 ;
			32'h00100f5c : data_o = 32'h06b3ffc8 ;
			32'h00100f60 : data_o = 32'h079340e6 ;
			32'h00100f64 : data_o = 32'hc8630200 ;
			32'h00100f68 : data_o = 32'h86ae06d7 ;
			32'h00100f6c : data_o = 32'h716387ba ;
			32'h00100f70 : data_o = 32'ha80302c7 ;
			32'h00100f74 : data_o = 32'h07910006 ;
			32'h00100f78 : data_o = 32'hae230691 ;
			32'h00100f7c : data_o = 32'heae3ff07 ;
			32'h00100f80 : data_o = 32'h0793fec7 ;
			32'h00100f84 : data_o = 32'h8f99fff6 ;
			32'h00100f88 : data_o = 32'h07919bf1 ;
			32'h00100f8c : data_o = 32'h95be973e ;
			32'h00100f90 : data_o = 32'h01176663 ;
			32'h00100f94 : data_o = 32'h872a8082 ;
			32'h00100f98 : data_o = 32'h03157e63 ;
			32'h00100f9c : data_o = 32'h0005c783 ;
			32'h00100fa0 : data_o = 32'h05850705 ;
			32'h00100fa4 : data_o = 32'hfef70fa3 ;
			32'h00100fa8 : data_o = 32'hfee89ae3 ;
			32'h00100fac : data_o = 32'hc6838082 ;
			32'h00100fb0 : data_o = 32'h07050005 ;
			32'h00100fb4 : data_o = 32'h00377793 ;
			32'h00100fb8 : data_o = 32'hfed70fa3 ;
			32'h00100fbc : data_o = 32'hdfd10585 ;
			32'h00100fc0 : data_o = 32'h0005c683 ;
			32'h00100fc4 : data_o = 32'h77930705 ;
			32'h00100fc8 : data_o = 32'h0fa30037 ;
			32'h00100fcc : data_o = 32'h0585fed7 ;
			32'h00100fd0 : data_o = 32'hb761fff9 ;
			32'h00100fd4 : data_o = 32'h11418082 ;
			32'h00100fd8 : data_o = 32'h0413c622 ;
			32'h00100fdc : data_o = 32'ha3830200 ;
			32'h00100fe0 : data_o = 32'ha2830005 ;
			32'h00100fe4 : data_o = 32'haf830045 ;
			32'h00100fe8 : data_o = 32'haf030085 ;
			32'h00100fec : data_o = 32'hae8300c5 ;
			32'h00100ff0 : data_o = 32'hae030105 ;
			32'h00100ff4 : data_o = 32'ha3030145 ;
			32'h00100ff8 : data_o = 32'ha8030185 ;
			32'h00100ffc : data_o = 32'h519401c5 ;
			32'h00101000 : data_o = 32'h02470713 ;
			32'h00101004 : data_o = 32'h40e607b3 ;
			32'h00101008 : data_o = 32'hfc772e23 ;
			32'h0010100c : data_o = 32'hfe572023 ;
			32'h00101010 : data_o = 32'hfff72223 ;
			32'h00101014 : data_o = 32'hffe72423 ;
			32'h00101018 : data_o = 32'hffd72623 ;
			32'h0010101c : data_o = 32'hffc72823 ;
			32'h00101020 : data_o = 32'hfe672a23 ;
			32'h00101024 : data_o = 32'hff072c23 ;
			32'h00101028 : data_o = 32'hfed72e23 ;
			32'h0010102c : data_o = 32'h02458593 ;
			32'h00101030 : data_o = 32'hfaf447e3 ;
			32'h00101034 : data_o = 32'h87ba86ae ;
			32'h00101038 : data_o = 32'h02c77163 ;
			32'h0010103c : data_o = 32'h0006a803 ;
			32'h00101040 : data_o = 32'h06910791 ;
			32'h00101044 : data_o = 32'hff07ae23 ;
			32'h00101048 : data_o = 32'hfec7eae3 ;
			32'h0010104c : data_o = 32'hfff60793 ;
			32'h00101050 : data_o = 32'h9bf18f99 ;
			32'h00101054 : data_o = 32'h973e0791 ;
			32'h00101058 : data_o = 32'h656395be ;
			32'h0010105c : data_o = 32'h44320117 ;
			32'h00101060 : data_o = 32'h80820141 ;
			32'h00101064 : data_o = 32'h0005c783 ;
			32'h00101068 : data_o = 32'h05850705 ;
			32'h0010106c : data_o = 32'hfef70fa3 ;
			32'h00101070 : data_o = 32'hfee887e3 ;
			32'h00101074 : data_o = 32'h0005c783 ;
			32'h00101078 : data_o = 32'h05850705 ;
			32'h0010107c : data_o = 32'hfef70fa3 ;
			32'h00101080 : data_o = 32'hfee892e3 ;
			32'h00101084 : data_o = 32'h0000bfe9 ;
			32'h00101088 : data_o = 32'he2de6f8d ;
			32'h0010108c : data_o = 32'h13880867 ;
			32'h00101090 : data_o = 32'h18af39e2 ;
			32'h00101094 : data_o = 32'hbc96e83f ;
			32'h00101098 : data_o = 32'he1e32beb ;
			32'h0010109c : data_o = 32'h3fd39163 ;
			32'h001010a0 : data_o = 32'hb82c818d ;
			32'h001010a4 : data_o = 32'h6845831c ;
			32'h001010a8 : data_o = 32'hdfe16d8e ;
			32'h001010ac : data_o = 32'h34783672 ;
			32'h001010b0 : data_o = 32'h1459e1f5 ;
			32'h001010b4 : data_o = 32'h456cd04d ;
			32'h001010b8 : data_o = 32'hd71e1fed ;
			32'h001010bc : data_o = 32'hf9cf77f1 ;
			32'h001010c0 : data_o = 32'h2c454c79 ;
			32'h001010c4 : data_o = 32'h76245b41 ;
			32'h001010c8 : data_o = 32'h072e47c9 ;
			32'h001010cc : data_o = 32'h1ce0b25c ;
			32'h001010d0 : data_o = 32'haf674757 ;
			32'h001010d4 : data_o = 32'h6d8d34cd ;
			32'h001010d8 : data_o = 32'h6e6c06b8 ;
			32'h001010dc : data_o = 32'h4431de61 ;
			32'h001010e0 : data_o = 32'he11ea286 ;
			32'h001010e4 : data_o = 32'hba2ef9ef ;
			32'h001010e8 : data_o = 32'hc36e84d9 ;
			32'h001010ec : data_o = 32'h387a1b10 ;
			32'h001010f0 : data_o = 32'h4db297c0 ;
			32'h001010f4 : data_o = 32'h431561cd ;
			32'h001010f8 : data_o = 32'hf7d817c2 ;
			32'h001010fc : data_o = 32'h0a394865 ;
			32'h00101100 : data_o = 32'h51d62a56 ;
			32'h00101104 : data_o = 32'hed72c725 ;
			32'h00101108 : data_o = 32'ha3e9e02e ;
			32'h0010110c : data_o = 32'hbb97ce6e ;
			32'h00101110 : data_o = 32'hc9372a22 ;
			32'h00101114 : data_o = 32'hc4d80cc4 ;
			32'h00101118 : data_o = 32'h39500671 ;
			32'h0010111c : data_o = 32'h6e12fa94 ;
			32'h00101120 : data_o = 32'h2ff6b8ed ;
			32'h00101124 : data_o = 32'ha625a7e5 ;
			32'h00101128 : data_o = 32'hffef2b46 ;
			32'h0010112c : data_o = 32'h27109969 ;
			32'h00101130 : data_o = 32'hb93ffc4a ;
			32'h00101134 : data_o = 32'h7725c985 ;
			32'h00101138 : data_o = 32'hd1c1f323 ;
			32'h0010113c : data_o = 32'h0e63e18f ;
			32'h00101140 : data_o = 32'he5a41796 ;
			32'h00101144 : data_o = 32'h20ba9d2b ;
			32'h00101148 : data_o = 32'hf290d99d ;
			32'h0010114c : data_o = 32'h3e4e945c ;
			32'h00101150 : data_o = 32'hf210cd15 ;
			32'h00101154 : data_o = 32'hf7b581f2 ;
			32'h00101158 : data_o = 32'h10d9624a ;
			32'h0010115c : data_o = 32'h34770359 ;
			32'h00101160 : data_o = 32'ha7f31e1f ;
			32'h00101164 : data_o = 32'ha621c285 ;
			32'h00101168 : data_o = 32'h4eb0c2c7 ;
			32'h0010116c : data_o = 32'h8fadfe18 ;
			32'h00101170 : data_o = 32'h3e389952 ;
			32'h00101174 : data_o = 32'h05d62f12 ;
			32'h00101178 : data_o = 32'h2264e879 ;
			32'h0010117c : data_o = 32'hd5909c4d ;
			32'h00101180 : data_o = 32'hdffd9cc1 ;
			32'h00101184 : data_o = 32'h25ed3e41 ;
			32'h00101188 : data_o = 32'hfd2987c2 ;
			32'h0010118c : data_o = 32'hc3e7739f ;
			32'h00101190 : data_o = 32'hc1402124 ;
			32'h00101194 : data_o = 32'hde5719b5 ;
			32'h00101198 : data_o = 32'he0191311 ;
			32'h0010119c : data_o = 32'h67a273a2 ;
			32'h001011a0 : data_o = 32'h362da406 ;
			32'h001011a4 : data_o = 32'h8e2fa366 ;
			32'h001011a8 : data_o = 32'hc06d9184 ;
			32'h001011ac : data_o = 32'hca6c4a75 ;
			32'h001011b0 : data_o = 32'h79567da3 ;
			32'h001011b4 : data_o = 32'h3cca7486 ;
			32'h001011b8 : data_o = 32'h8f7d6e1f ;
			32'h001011bc : data_o = 32'haaac1d55 ;
			32'h001011c0 : data_o = 32'hb39ebc43 ;
			32'h001011c4 : data_o = 32'hf17fb474 ;
			32'h001011c8 : data_o = 32'hfa6fa8ca ;
			32'h001011cc : data_o = 32'h79cb4b80 ;
			32'h001011d0 : data_o = 32'hbf12ba96 ;
			32'h001011d4 : data_o = 32'h514fbd7d ;
			32'h001011d8 : data_o = 32'h0b6b45b1 ;
			32'h001011dc : data_o = 32'h609b967b ;
			32'h001011e0 : data_o = 32'hc8b5fd54 ;
			32'h001011e4 : data_o = 32'hf9341c56 ;
			32'h001011e8 : data_o = 32'hea7b657d ;
			32'h001011ec : data_o = 32'h9fb10d4c ;
			32'h001011f0 : data_o = 32'h9a9f4f6d ;
			32'h001011f4 : data_o = 32'hab8f81c6 ;
			32'h001011f8 : data_o = 32'h27b5f004 ;
			32'h001011fc : data_o = 32'ha5daad14 ;
			32'h00101200 : data_o = 32'h4c56f386 ;
			32'h00101204 : data_o = 32'h481a4830 ;
			32'h00101208 : data_o = 32'hce3dee17 ;
			32'h0010120c : data_o = 32'he5d1ad2f ;
			32'h00101210 : data_o = 32'h277041c5 ;
			32'h00101214 : data_o = 32'hbd36865d ;
			32'h00101218 : data_o = 32'h9c7f6486 ;
			32'h0010121c : data_o = 32'h928a3a7f ;
			32'h00101220 : data_o = 32'h84fbe4e1 ;
			32'h00101224 : data_o = 32'habe83be0 ;
			32'h00101228 : data_o = 32'h0202ea99 ;
			32'h0010122c : data_o = 32'hc0fc1e75 ;
			32'h00101230 : data_o = 32'hf7495dc1 ;
			32'h00101234 : data_o = 32'hbe0d9b9c ;
			32'h00101238 : data_o = 32'h65151d5d ;
			32'h0010123c : data_o = 32'h47deeb16 ;
			32'h00101240 : data_o = 32'h15b9e4ae ;
			32'h00101244 : data_o = 32'hb51d48d3 ;
			32'h00101248 : data_o = 32'h8e139b5b ;
			32'h0010124c : data_o = 32'hddbd4422 ;
			32'h00101250 : data_o = 32'h091ff5e0 ;
			32'h00101254 : data_o = 32'h53de9c72 ;
			32'h00101258 : data_o = 32'h9773cfda ;
			32'h0010125c : data_o = 32'h15d93ec5 ;
			32'h00101260 : data_o = 32'h7159361c ;
			32'h00101264 : data_o = 32'h753d49ef ;
			32'h00101268 : data_o = 32'hb37c5e6c ;
			32'h0010126c : data_o = 32'h0e82c85d ;
			32'h00101270 : data_o = 32'h13aad8ec ;
			32'h00101274 : data_o = 32'h33e6ddb7 ;
			32'h00101278 : data_o = 32'h2d9e6e03 ;
			32'h0010127c : data_o = 32'hb3d2855f ;
			32'h00101280 : data_o = 32'h99b46431 ;
			32'h00101284 : data_o = 32'h37b49fd2 ;
			32'h00101288 : data_o = 32'h76504d9e ;
			32'h0010128c : data_o = 32'h8fa390aa ;
			32'h00101290 : data_o = 32'hf5047742 ;
			32'h00101294 : data_o = 32'h40bf7c79 ;
			32'h00101298 : data_o = 32'hd705e1c6 ;
			32'h0010129c : data_o = 32'h4dbd96e5 ;
			32'h001012a0 : data_o = 32'h4863ead2 ;
			32'h001012a4 : data_o = 32'h94d7e57f ;
			32'h001012a8 : data_o = 32'h5c9997ab ;
			32'h001012ac : data_o = 32'h296adf06 ;
			32'h001012b0 : data_o = 32'h60ec814c ;
			32'h001012b4 : data_o = 32'he7e13a0a ;
			32'h001012b8 : data_o = 32'h9f96ae87 ;
			32'h001012bc : data_o = 32'h5899d4f7 ;
			32'h001012c0 : data_o = 32'h6cad386b ;
			32'h001012c4 : data_o = 32'h66df6fe2 ;
			32'h001012c8 : data_o = 32'h657ff310 ;
			32'h001012cc : data_o = 32'h79929904 ;
			32'h001012d0 : data_o = 32'h7756c292 ;
			32'h001012d4 : data_o = 32'h6c9c2301 ;
			32'h001012d8 : data_o = 32'haf282fbe ;
			32'h001012dc : data_o = 32'h67cebd30 ;
			32'h001012e0 : data_o = 32'h65e33775 ;
			32'h001012e4 : data_o = 32'h8fb0a281 ;
			32'h001012e8 : data_o = 32'h414d7fc9 ;
			32'h001012ec : data_o = 32'h9bff939a ;
			32'h001012f0 : data_o = 32'hf295af9c ;
			32'h001012f4 : data_o = 32'h3e5aea74 ;
			32'h001012f8 : data_o = 32'h6139d318 ;
			32'h001012fc : data_o = 32'h1d550395 ;
			32'h00101300 : data_o = 32'ha4a069e1 ;
			32'h00101304 : data_o = 32'he3f0ef5c ;
			32'h00101308 : data_o = 32'h040c854d ;
			32'h0010130c : data_o = 32'h988bdc62 ;
			32'h00101310 : data_o = 32'hdebd9e9c ;
			32'h00101314 : data_o = 32'hb3493868 ;
			32'h00101318 : data_o = 32'h787b5bc4 ;
			32'h0010131c : data_o = 32'hbcd85312 ;
			32'h00101320 : data_o = 32'hd0328121 ;
			32'h00101324 : data_o = 32'h0b04b427 ;
			32'h00101328 : data_o = 32'h8c4e468c ;
			32'h0010132c : data_o = 32'h1a1e0630 ;
			32'h00101330 : data_o = 32'h97848520 ;
			32'h00101334 : data_o = 32'h4cf7e4bc ;
			32'h00101338 : data_o = 32'hb338c8ab ;
			32'h0010133c : data_o = 32'habde3dd6 ;
			32'h00101340 : data_o = 32'h2a75cf62 ;
			32'h00101344 : data_o = 32'hb3398c9d ;
			32'h00101348 : data_o = 32'h19f220dd ;
			32'h0010134c : data_o = 32'hf19e096c ;
			32'h00101350 : data_o = 32'hc9a50292 ;
			32'h00101354 : data_o = 32'h69f5d974 ;
			32'h00101358 : data_o = 32'hf2e8104c ;
			32'h0010135c : data_o = 32'h7123eae4 ;
			32'h00101360 : data_o = 32'hce7d32ed ;
			32'h00101364 : data_o = 32'h9b1cee5b ;
			32'h00101368 : data_o = 32'hd262d97c ;
			32'h0010136c : data_o = 32'h77472e2c ;
			32'h00101370 : data_o = 32'h6bc6d945 ;
			32'h00101374 : data_o = 32'h92d4246a ;
			32'h00101378 : data_o = 32'hb515e17d ;
			32'h0010137c : data_o = 32'hc3d91256 ;
			32'h00101380 : data_o = 32'hc9474ad6 ;
			32'h00101384 : data_o = 32'hd2c01c04 ;
			32'h00101388 : data_o = 32'h0fb62692 ;
			32'h0010138c : data_o = 32'h63f79fcd ;
			32'h00101390 : data_o = 32'hebb21e00 ;
			32'h00101394 : data_o = 32'h5400bb82 ;
			32'h00101398 : data_o = 32'ha5153d38 ;
			32'h0010139c : data_o = 32'hde573ca7 ;
			32'h001013a0 : data_o = 32'h1f120428 ;
			32'h001013a4 : data_o = 32'hcd00473f ;
			32'h001013a8 : data_o = 32'h4b49d242 ;
			32'h001013ac : data_o = 32'ha59cb88c ;
			32'h001013b0 : data_o = 32'h8f39f6b0 ;
			32'h001013b4 : data_o = 32'h21061ff5 ;
			32'h001013b8 : data_o = 32'hda0320c4 ;
			32'h001013bc : data_o = 32'hd74eb543 ;
			32'h001013c0 : data_o = 32'h370b5f33 ;
			32'h001013c4 : data_o = 32'h2731248d ;
			32'h001013c8 : data_o = 32'had860b93 ;
			32'h001013cc : data_o = 32'h572c21d5 ;
			32'h001013d0 : data_o = 32'h2ed33c79 ;
			32'h001013d4 : data_o = 32'ha24d2a17 ;
			32'h001013d8 : data_o = 32'h617074a7 ;
			32'h001013dc : data_o = 32'he2fe149f ;
			32'h001013e0 : data_o = 32'h7acdbc28 ;
			32'h001013e4 : data_o = 32'h1ce6557a ;
			32'h001013e8 : data_o = 32'h8b75a5c1 ;
			32'h001013ec : data_o = 32'hae515a4c ;
			32'h001013f0 : data_o = 32'h85b5130a ;
			32'h001013f4 : data_o = 32'h2810fc90 ;
			32'h001013f8 : data_o = 32'heac0620c ;
			32'h001013fc : data_o = 32'h68dc4430 ;
			32'h00101400 : data_o = 32'h2e13d678 ;
			32'h00101404 : data_o = 32'hf28fcea6 ;
			32'h00101408 : data_o = 32'h10ec1d20 ;
			32'h0010140c : data_o = 32'ha7e41f8a ;
			32'h00101410 : data_o = 32'h8e8db786 ;
			32'h00101414 : data_o = 32'he8ada5d1 ;
			32'h00101418 : data_o = 32'h34ae2b5a ;
			32'h0010141c : data_o = 32'h64339042 ;
			32'h00101420 : data_o = 32'h5d999bd1 ;
			32'h00101424 : data_o = 32'hff739ce7 ;
			32'h00101428 : data_o = 32'h96f523ee ;
			32'h0010142c : data_o = 32'h34b4202b ;
			32'h00101430 : data_o = 32'h276d5fa1 ;
			32'h00101434 : data_o = 32'hf9fba74e ;
			32'h00101438 : data_o = 32'h43121cc3 ;
			32'h0010143c : data_o = 32'h63467def ;
			32'h00101440 : data_o = 32'hf709b61e ;
			32'h00101444 : data_o = 32'h0ffdf0be ;
			32'h00101448 : data_o = 32'hec10e79b ;
			32'h0010144c : data_o = 32'h741bc4a6 ;
			32'h00101450 : data_o = 32'h37a59906 ;
			32'h00101454 : data_o = 32'h377f9492 ;
			32'h00101458 : data_o = 32'h55f970d1 ;
			32'h0010145c : data_o = 32'hba8a32d7 ;
			32'h00101460 : data_o = 32'ha3881619 ;
			32'h00101464 : data_o = 32'hddb69378 ;
			32'h00101468 : data_o = 32'h629b235f ;
			32'h0010146c : data_o = 32'h67a9cb91 ;
			32'h00101470 : data_o = 32'h3732582a ;
			32'h00101474 : data_o = 32'h639dd874 ;
			32'h00101478 : data_o = 32'h054a20f1 ;
			32'h0010147c : data_o = 32'h5ab9f30a ;
			32'h00101480 : data_o = 32'hff158acf ;
			32'h00101484 : data_o = 32'h16aeaa59 ;
			32'h00101488 : data_o = 32'h813c716c ;
			32'h0010148c : data_o = 32'hb04af7c7 ;
			32'h00101490 : data_o = 32'h9cd4f1ec ;
			32'h00101494 : data_o = 32'h0b41f4d5 ;
			32'h00101498 : data_o = 32'h6d33a13f ;
			32'h0010149c : data_o = 32'hbbd0a9e1 ;
			32'h001014a0 : data_o = 32'hb4425ab2 ;
			32'h001014a4 : data_o = 32'hb1f8885b ;
			32'h001014a8 : data_o = 32'h917f6d9c ;
			32'h001014ac : data_o = 32'hb14b517a ;
			32'h001014b0 : data_o = 32'hec7afd4b ;
			32'h001014b4 : data_o = 32'hd5179f0a ;
			32'h001014b8 : data_o = 32'h73824909 ;
			32'h001014bc : data_o = 32'h9bbe37fb ;
			32'h001014c0 : data_o = 32'ha2c77e00 ;
			32'h001014c4 : data_o = 32'hcc514c90 ;
			32'h001014c8 : data_o = 32'hd689d0da ;
			32'h001014cc : data_o = 32'h5af9fe14 ;
			32'h001014d0 : data_o = 32'he88c9005 ;
			32'h001014d4 : data_o = 32'hbe50d5a9 ;
			32'h001014d8 : data_o = 32'h1f5bd890 ;
			32'h001014dc : data_o = 32'h0e9e3b7a ;
			32'h001014e0 : data_o = 32'h55126e06 ;
			32'h001014e4 : data_o = 32'hbf104e35 ;
			32'h001014e8 : data_o = 32'h32958900 ;
			32'h001014ec : data_o = 32'h35f201c1 ;
			32'h001014f0 : data_o = 32'hf23384d6 ;
			32'h001014f4 : data_o = 32'h1766e24d ;
			32'h001014f8 : data_o = 32'hba4ebbf5 ;
			32'h001014fc : data_o = 32'ha125028d ;
			32'h00101500 : data_o = 32'hb075c458 ;
			32'h00101504 : data_o = 32'h7f9f93bf ;
			32'h00101508 : data_o = 32'h6dad577f ;
			32'h0010150c : data_o = 32'h5daeb54d ;
			32'h00101510 : data_o = 32'h8796698e ;
			32'h00101514 : data_o = 32'h07ffc6dc ;
			32'h00101518 : data_o = 32'hf1d889a8 ;
			32'h0010151c : data_o = 32'h1303dead ;
			32'h00101520 : data_o = 32'h71c3161f ;
			32'h00101524 : data_o = 32'h45db58ab ;
			32'h00101528 : data_o = 32'hd8a69ad1 ;
			32'h0010152c : data_o = 32'h0270b695 ;
			32'h00101530 : data_o = 32'h09a09743 ;
			32'h00101534 : data_o = 32'h4e692812 ;
			32'h00101538 : data_o = 32'h6cf32b26 ;
			32'h0010153c : data_o = 32'h21457d36 ;
			32'h00101540 : data_o = 32'h7ff2e0c2 ;
			32'h00101544 : data_o = 32'h222a4907 ;
			32'h00101548 : data_o = 32'hab8aac79 ;
			32'h0010154c : data_o = 32'h639dec8f ;
			32'h00101550 : data_o = 32'hd99c4eba ;
			32'h00101554 : data_o = 32'haf688035 ;
			32'h00101558 : data_o = 32'hffc4d5c2 ;
			32'h0010155c : data_o = 32'h8eb5f536 ;
			32'h00101560 : data_o = 32'ha883c311 ;
			32'h00101564 : data_o = 32'h1dc5d32d ;
			32'h00101568 : data_o = 32'hc1ff2501 ;
			32'h0010156c : data_o = 32'hd12db6c0 ;
			32'h00101570 : data_o = 32'hc204953d ;
			32'h00101574 : data_o = 32'h4f8c3c87 ;
			32'h00101578 : data_o = 32'h5ace9a39 ;
			32'h0010157c : data_o = 32'hed822dce ;
			32'h00101580 : data_o = 32'hfd4f56b4 ;
			32'h00101584 : data_o = 32'h53c91684 ;
			32'h00101588 : data_o = 32'h3e125fa3 ;
			32'h0010158c : data_o = 32'ha8bee20b ;
			32'h00101590 : data_o = 32'heaf7a5ee ;
			32'h00101594 : data_o = 32'h003e44db ;
			32'h00101598 : data_o = 32'hd640f373 ;
			32'h0010159c : data_o = 32'h796f2058 ;
			32'h001015a0 : data_o = 32'h5d0564a8 ;
			32'h001015a4 : data_o = 32'h7320373f ;
			32'h001015a8 : data_o = 32'h91564186 ;
			32'h001015ac : data_o = 32'h3933e450 ;
			32'h001015b0 : data_o = 32'h1dabc6a8 ;
			32'h001015b4 : data_o = 32'hd5a52fae ;
			32'h001015b8 : data_o = 32'h4182dbe3 ;
			32'h001015bc : data_o = 32'hde514117 ;
			32'h001015c0 : data_o = 32'h620254c3 ;
			32'h001015c4 : data_o = 32'h131f73d9 ;
			32'h001015c8 : data_o = 32'h9ea14e99 ;
			32'h001015cc : data_o = 32'h84cfad5d ;
			32'h001015d0 : data_o = 32'hacc2f8a2 ;
			32'h001015d4 : data_o = 32'h834246ee ;
			32'h001015d8 : data_o = 32'h2970d5bf ;
			32'h001015dc : data_o = 32'h2ff6a9a0 ;
			32'h001015e0 : data_o = 32'h3c6c66ab ;
			32'h001015e4 : data_o = 32'hd73904cc ;
			32'h001015e8 : data_o = 32'ha1f6f687 ;
			32'h001015ec : data_o = 32'hfce09402 ;
			32'h001015f0 : data_o = 32'hfe9b5b6b ;
			32'h001015f4 : data_o = 32'h6d278d37 ;
			32'h001015f8 : data_o = 32'h4b1246b0 ;
			32'h001015fc : data_o = 32'h2034e2bf ;
			32'h00101600 : data_o = 32'h0dd80b57 ;
			32'h00101604 : data_o = 32'hb3257cf2 ;
			32'h00101608 : data_o = 32'hf4a6ec31 ;
			32'h0010160c : data_o = 32'h0d107446 ;
			32'h00101610 : data_o = 32'h3f762ce6 ;
			32'h00101614 : data_o = 32'h2279802c ;
			32'h00101618 : data_o = 32'h7cc84b08 ;
			32'h0010161c : data_o = 32'hadb6d8ff ;
			32'h00101620 : data_o = 32'ha7848d35 ;
			32'h00101624 : data_o = 32'hc70952fa ;
			32'h00101628 : data_o = 32'hee8aff4a ;
			32'h0010162c : data_o = 32'hf27a19e3 ;
			32'h00101630 : data_o = 32'hb07a1918 ;
			32'h00101634 : data_o = 32'hca3aada1 ;
			32'h00101638 : data_o = 32'hebfbba70 ;
			32'h0010163c : data_o = 32'h412fe212 ;
			32'h00101640 : data_o = 32'hfb8d725c ;
			32'h00101644 : data_o = 32'h7302b5af ;
			32'h00101648 : data_o = 32'hf5b7911c ;
			32'h0010164c : data_o = 32'hc527e37b ;
			32'h00101650 : data_o = 32'h99fb1352 ;
			32'h00101654 : data_o = 32'h5d471e3d ;
			32'h00101658 : data_o = 32'haea1a3ac ;
			32'h0010165c : data_o = 32'h69c696d5 ;
			32'h00101660 : data_o = 32'h55d884eb ;
			32'h00101664 : data_o = 32'h1c912784 ;
			32'h00101668 : data_o = 32'hb475cd57 ;
			32'h0010166c : data_o = 32'h1bceff61 ;
			32'h00101670 : data_o = 32'h897e8a16 ;
			32'h00101674 : data_o = 32'hd0e1455a ;
			32'h00101678 : data_o = 32'hf738e194 ;
			32'h0010167c : data_o = 32'h5f5f866b ;
			32'h00101680 : data_o = 32'hb80d0242 ;
			32'h00101684 : data_o = 32'h92b9b8a9 ;
			32'h00101688 : data_o = 32'h9c8c993f ;
			32'h0010168c : data_o = 32'hcc4e2f2c ;
			32'h00101690 : data_o = 32'h8f28ff5a ;
			32'h00101694 : data_o = 32'hfe26b5ed ;
			32'h00101698 : data_o = 32'h6d9c130b ;
			32'h0010169c : data_o = 32'hf975526d ;
			32'h001016a0 : data_o = 32'h8e087e22 ;
			32'h001016a4 : data_o = 32'h0c39effa ;
			32'h001016a8 : data_o = 32'h495ff12b ;
			32'h001016ac : data_o = 32'h9506cb98 ;
			32'h001016b0 : data_o = 32'h75d3ee52 ;
			32'h001016b4 : data_o = 32'h8a414622 ;
			32'h001016b8 : data_o = 32'h7d34a985 ;
			32'h001016bc : data_o = 32'h64f2d84c ;
			32'h001016c0 : data_o = 32'h345e5693 ;
			32'h001016c4 : data_o = 32'h8947fe45 ;
			32'h001016c8 : data_o = 32'h08751946 ;
			32'h001016cc : data_o = 32'heaf1c6d0 ;
			32'h001016d0 : data_o = 32'h3ac777d8 ;
			32'h001016d4 : data_o = 32'h7311b459 ;
			32'h001016d8 : data_o = 32'h4499a187 ;
			32'h001016dc : data_o = 32'hccff9451 ;
			32'h001016e0 : data_o = 32'h1c29e0d5 ;
			32'h001016e4 : data_o = 32'ha9f3a082 ;
			32'h001016e8 : data_o = 32'h9ee65720 ;
			32'h001016ec : data_o = 32'h92cf31c0 ;
			32'h001016f0 : data_o = 32'h8b3c69f4 ;
			32'h001016f4 : data_o = 32'h37410c9b ;
			32'h001016f8 : data_o = 32'hdd55018b ;
			32'h001016fc : data_o = 32'h98010bf6 ;
			32'h00101700 : data_o = 32'hcfb78838 ;
			32'h00101704 : data_o = 32'h587025e7 ;
			32'h00101708 : data_o = 32'ha93d4a23 ;
			32'h0010170c : data_o = 32'h216636e0 ;
			32'h00101710 : data_o = 32'h648c137a ;
			32'h00101714 : data_o = 32'h8cbdad57 ;
			32'h00101718 : data_o = 32'h5ca7e3ae ;
			32'h0010171c : data_o = 32'h8c118469 ;
			32'h00101720 : data_o = 32'hdacf7414 ;
			32'h00101724 : data_o = 32'hed8ff046 ;
			32'h00101728 : data_o = 32'h65976130 ;
			32'h0010172c : data_o = 32'h9b87966c ;
			32'h00101730 : data_o = 32'hb0cc6562 ;
			32'h00101734 : data_o = 32'hd64c3f39 ;
			32'h00101738 : data_o = 32'h8204a7f2 ;
			32'h0010173c : data_o = 32'hf3232b96 ;
			32'h00101740 : data_o = 32'h53afe6d0 ;
			32'h00101744 : data_o = 32'h9207e9ff ;
			32'h00101748 : data_o = 32'he28a6d3e ;
			32'h0010174c : data_o = 32'h2c967a3c ;
			32'h00101750 : data_o = 32'h9895bee1 ;
			32'h00101754 : data_o = 32'h4e31eecb ;
			32'h00101758 : data_o = 32'hc9129637 ;
			32'h0010175c : data_o = 32'h6af2048c ;
			32'h00101760 : data_o = 32'h03d02ddc ;
			32'h00101764 : data_o = 32'hc1d24387 ;
			32'h00101768 : data_o = 32'h6eb7391d ;
			32'h0010176c : data_o = 32'h576bfc8d ;
			32'h00101770 : data_o = 32'h8c8a9283 ;
			32'h00101774 : data_o = 32'h6a9bcc7a ;
			32'h00101778 : data_o = 32'hee6df2a0 ;
			32'h0010177c : data_o = 32'hfc054586 ;
			32'h00101780 : data_o = 32'h270b148c ;
			32'h00101784 : data_o = 32'h8eab0e30 ;
			32'h00101788 : data_o = 32'h8736face ;
			32'h0010178c : data_o = 32'hf1920353 ;
			32'h00101790 : data_o = 32'h0fbc8007 ;
			32'h00101794 : data_o = 32'h10c13e21 ;
			32'h00101798 : data_o = 32'h2692061d ;
			32'h0010179c : data_o = 32'h20730e6d ;
			32'h001017a0 : data_o = 32'h74fd194d ;
			32'h001017a4 : data_o = 32'h1e9aaf15 ;
			32'h001017a8 : data_o = 32'hf7d38c38 ;
			32'h001017ac : data_o = 32'h930e7d9b ;
			32'h001017b0 : data_o = 32'h1e73bdee ;
			32'h001017b4 : data_o = 32'hbff67e85 ;
			32'h001017b8 : data_o = 32'h22b0ce0e ;
			32'h001017bc : data_o = 32'h7575c9b2 ;
			32'h001017c0 : data_o = 32'hbbebcccc ;
			32'h001017c4 : data_o = 32'h46b0b28b ;
			32'h001017c8 : data_o = 32'h6008d540 ;
			32'h001017cc : data_o = 32'h7ca7f08d ;
			32'h001017d0 : data_o = 32'he25567b1 ;
			32'h001017d4 : data_o = 32'h79f9fed8 ;
			32'h001017d8 : data_o = 32'h827056d0 ;
			32'h001017dc : data_o = 32'h1abd103f ;
			32'h001017e0 : data_o = 32'h0dddbc64 ;
			32'h001017e4 : data_o = 32'hbd397276 ;
			32'h001017e8 : data_o = 32'h6ce4a3a3 ;
			32'h001017ec : data_o = 32'hf2b3c84b ;
			32'h001017f0 : data_o = 32'ha1fe3abe ;
			32'h001017f4 : data_o = 32'h29c7f7e9 ;
			32'h001017f8 : data_o = 32'hb2f91184 ;
			32'h001017fc : data_o = 32'hd2f14cbd ;
			32'h00101800 : data_o = 32'h1c8377f0 ;
			32'h00101804 : data_o = 32'h0244d8de ;
			32'h00101808 : data_o = 32'he043927d ;
			32'h0010180c : data_o = 32'h9e270462 ;
			32'h00101810 : data_o = 32'hae0d0184 ;
			32'h00101814 : data_o = 32'h30d33574 ;
			32'h00101818 : data_o = 32'hd1ea6358 ;
			32'h0010181c : data_o = 32'ha6fa9a74 ;
			32'h00101820 : data_o = 32'h3395a5f8 ;
			32'h00101824 : data_o = 32'h8e515d9c ;
			32'h00101828 : data_o = 32'h75217b81 ;
			32'h0010182c : data_o = 32'he9cbb804 ;
			32'h00101830 : data_o = 32'h675eedd5 ;
			32'h00101834 : data_o = 32'h71376a7b ;
			32'h00101838 : data_o = 32'h155f9f76 ;
			32'h0010183c : data_o = 32'h642c92a4 ;
			32'h00101840 : data_o = 32'hd2b29395 ;
			32'h00101844 : data_o = 32'hb1334016 ;
			32'h00101848 : data_o = 32'hb2e79a59 ;
			32'h0010184c : data_o = 32'hae717491 ;
			32'h00101850 : data_o = 32'h6a119861 ;
			32'h00101854 : data_o = 32'hd50fc061 ;
			32'h00101858 : data_o = 32'hed1b9bac ;
			32'h0010185c : data_o = 32'hebcd88c6 ;
			32'h00101860 : data_o = 32'ha6c0836a ;
			32'h00101864 : data_o = 32'h6fa28302 ;
			32'h00101868 : data_o = 32'hc59b4e61 ;
			32'h0010186c : data_o = 32'ha2e74e76 ;
			32'h00101870 : data_o = 32'had0f7213 ;
			32'h00101874 : data_o = 32'he9352df4 ;
			32'h00101878 : data_o = 32'h6edd5813 ;
			32'h0010187c : data_o = 32'hf85c9e7c ;
			32'h00101880 : data_o = 32'hac75f5ba ;
			32'h00101884 : data_o = 32'h06a0f35c ;
			32'h00101888 : data_o = 32'ha567805f ;
			32'h0010188c : data_o = 32'ha034571f ;
			32'h00101890 : data_o = 32'hd1718609 ;
			32'h00101894 : data_o = 32'h5aba658f ;
			32'h00101898 : data_o = 32'hcbd10168 ;
			32'h0010189c : data_o = 32'h271ecee5 ;
			32'h001018a0 : data_o = 32'h07afda6a ;
			32'h001018a4 : data_o = 32'h8bba88d2 ;
			32'h001018a8 : data_o = 32'ha534bcbc ;
			32'h001018ac : data_o = 32'h869d23f4 ;
			32'h001018b0 : data_o = 32'h2b296924 ;
			32'h001018b4 : data_o = 32'h95956895 ;
			32'h001018b8 : data_o = 32'h1ec973d4 ;
			32'h001018bc : data_o = 32'h05ed7418 ;
			32'h001018c0 : data_o = 32'h6403b37e ;
			32'h001018c4 : data_o = 32'h97b735c3 ;
			32'h001018c8 : data_o = 32'hc8ca0fdf ;
			32'h001018cc : data_o = 32'h8f066746 ;
			32'h001018d0 : data_o = 32'h21bb0044 ;
			32'h001018d4 : data_o = 32'hcc2c3526 ;
			32'h001018d8 : data_o = 32'hd279e5ed ;
			32'h001018dc : data_o = 32'h6ce92497 ;
			32'h001018e0 : data_o = 32'h2487b461 ;
			32'h001018e4 : data_o = 32'h6fd862bb ;
			32'h001018e8 : data_o = 32'hfdbbe865 ;
			32'h001018ec : data_o = 32'h6a519591 ;
			32'h001018f0 : data_o = 32'h23859157 ;
			32'h001018f4 : data_o = 32'hd92c5767 ;
			32'h001018f8 : data_o = 32'h2b3775c7 ;
			32'h001018fc : data_o = 32'h6c7c6717 ;
			32'h00101900 : data_o = 32'h406da1aa ;
			32'h00101904 : data_o = 32'h0e933f4b ;
			32'h00101908 : data_o = 32'h76cf40c9 ;
			32'h0010190c : data_o = 32'h5db3e454 ;
			32'h00101910 : data_o = 32'hcfcf8bc3 ;
			32'h00101914 : data_o = 32'ha98d7a94 ;
			32'h00101918 : data_o = 32'h0383c88c ;
			32'h0010191c : data_o = 32'hc7c8f8bc ;
			32'h00101920 : data_o = 32'he7b38b96 ;
			32'h00101924 : data_o = 32'hdfa38cbd ;
			32'h00101928 : data_o = 32'ha936392f ;
			32'h0010192c : data_o = 32'hba79db0c ;
			32'h00101930 : data_o = 32'h6f2c129d ;
			32'h00101934 : data_o = 32'h4a16f9d3 ;
			32'h00101938 : data_o = 32'hf7178252 ;
			32'h0010193c : data_o = 32'h74536a00 ;
			32'h00101940 : data_o = 32'h7d3291c1 ;
			32'h00101944 : data_o = 32'hf43db453 ;
			32'h00101948 : data_o = 32'h16fef98f ;
			32'h0010194c : data_o = 32'hc566d1de ;
			32'h00101950 : data_o = 32'hc3e9f2bd ;
			32'h00101954 : data_o = 32'h474fd263 ;
			32'h00101958 : data_o = 32'h30ec68ba ;
			32'h0010195c : data_o = 32'h957f93e5 ;
			32'h00101960 : data_o = 32'h427c5920 ;
			32'h00101964 : data_o = 32'ha1020de3 ;
			32'h00101968 : data_o = 32'h6794154c ;
			32'h0010196c : data_o = 32'h391ce65e ;
			32'h00101970 : data_o = 32'h294023aa ;
			32'h00101974 : data_o = 32'hb04859e2 ;
			32'h00101978 : data_o = 32'h62b8c612 ;
			32'h0010197c : data_o = 32'hcbe75321 ;
			32'h00101980 : data_o = 32'h2f3dbfc0 ;
			32'h00101984 : data_o = 32'h809765e5 ;
			32'h00101988 : data_o = 32'he230499a ;
			32'h0010198c : data_o = 32'h2e908990 ;
			32'h00101990 : data_o = 32'hf62e283c ;
			32'h00101994 : data_o = 32'hb37ebf78 ;
			32'h00101998 : data_o = 32'hc8ba6c07 ;
			32'h0010199c : data_o = 32'had97b95b ;
			32'h001019a0 : data_o = 32'h6287edce ;
			32'h001019a4 : data_o = 32'h7e02494a ;
			32'h001019a8 : data_o = 32'h8902ecd4 ;
			32'h001019ac : data_o = 32'hb468bb64 ;
			32'h001019b0 : data_o = 32'hc00c972f ;
			32'h001019b4 : data_o = 32'h930d6449 ;
			32'h001019b8 : data_o = 32'h78aa7811 ;
			32'h001019bc : data_o = 32'h2f425e22 ;
			32'h001019c0 : data_o = 32'h8d11e6b2 ;
			32'h001019c4 : data_o = 32'h0d9dc11e ;
			32'h001019c8 : data_o = 32'h08428d9d ;
			32'h001019cc : data_o = 32'h9f8080bb ;
			32'h001019d0 : data_o = 32'h37ce2792 ;
			32'h001019d4 : data_o = 32'h7a45119d ;
			32'h001019d8 : data_o = 32'hef92d137 ;
			32'h001019dc : data_o = 32'h50f8eb0c ;
			32'h001019e0 : data_o = 32'ha30dca74 ;
			32'h001019e4 : data_o = 32'h654390a5 ;
			32'h001019e8 : data_o = 32'h1dd07635 ;
			32'h001019ec : data_o = 32'h6c2f1de2 ;
			32'h001019f0 : data_o = 32'h0509d1ef ;
			32'h001019f4 : data_o = 32'h05c58e95 ;
			32'h001019f8 : data_o = 32'h04d88656 ;
			32'h001019fc : data_o = 32'haa9930e8 ;
			32'h00101a00 : data_o = 32'hf7394917 ;
			32'h00101a04 : data_o = 32'hfbf917ce ;
			32'h00101a08 : data_o = 32'hdeae4223 ;
			32'h00101a0c : data_o = 32'h5582aa2d ;
			32'h00101a10 : data_o = 32'h4d7ed00b ;
			32'h00101a14 : data_o = 32'h2d8e2778 ;
			32'h00101a18 : data_o = 32'h6746dc03 ;
			32'h00101a1c : data_o = 32'h91884bd4 ;
			32'h00101a20 : data_o = 32'h2c0565aa ;
			32'h00101a24 : data_o = 32'h3fc0a893 ;
			32'h00101a28 : data_o = 32'h4f0191cf ;
			32'h00101a2c : data_o = 32'he370c2b9 ;
			32'h00101a30 : data_o = 32'h97fff858 ;
			32'h00101a34 : data_o = 32'h7ce35f48 ;
			32'h00101a38 : data_o = 32'h62f021b4 ;
			32'h00101a3c : data_o = 32'h0adab08b ;
			32'h00101a40 : data_o = 32'h2fce77d9 ;
			32'h00101a44 : data_o = 32'hbabee02d ;
			32'h00101a48 : data_o = 32'hd23f6e19 ;
			32'h00101a4c : data_o = 32'h1e13d9f2 ;
			32'h00101a50 : data_o = 32'h276b68fb ;
			32'h00101a54 : data_o = 32'hff38f1de ;
			32'h00101a58 : data_o = 32'h342ada8a ;
			32'h00101a5c : data_o = 32'he311327b ;
			32'h00101a60 : data_o = 32'h6275062e ;
			32'h00101a64 : data_o = 32'h4dfc1299 ;
			32'h00101a68 : data_o = 32'h818afb52 ;
			32'h00101a6c : data_o = 32'h51a69489 ;
			32'h00101a70 : data_o = 32'heb277cbd ;
			32'h00101a74 : data_o = 32'hee240582 ;
			32'h00101a78 : data_o = 32'hfefaece1 ;
			32'h00101a7c : data_o = 32'h3b3f2a4b ;
			32'h00101a80 : data_o = 32'h4bf46921 ;
			32'h00101a84 : data_o = 32'hc7894bab ;
			32'h00101a88 : data_o = 32'h9388fd41 ;
			32'h00101a8c : data_o = 32'h26f289c3 ;
			32'h00101a90 : data_o = 32'h01666b90 ;
			32'h00101a94 : data_o = 32'hb73a9f5d ;
			32'h00101a98 : data_o = 32'h53cd8b41 ;
			32'h00101a9c : data_o = 32'hbae0d7bb ;
			32'h00101aa0 : data_o = 32'hc9e53c28 ;
			32'h00101aa4 : data_o = 32'hac9e955e ;
			32'h00101aa8 : data_o = 32'had43c6ed ;
			32'h00101aac : data_o = 32'h7854039b ;
			32'h00101ab0 : data_o = 32'h97267015 ;
			32'h00101ab4 : data_o = 32'h7c1d0dfc ;
			32'h00101ab8 : data_o = 32'hf399229f ;
			32'h00101abc : data_o = 32'h206fae2b ;
			32'h00101ac0 : data_o = 32'h4363165e ;
			32'h00101ac4 : data_o = 32'haac5ec36 ;
			32'h00101ac8 : data_o = 32'h92ebe375 ;
			32'h00101acc : data_o = 32'h227d4ef2 ;
			32'h00101ad0 : data_o = 32'hfac52b2c ;
			32'h00101ad4 : data_o = 32'hd6357443 ;
			32'h00101ad8 : data_o = 32'h8adbd977 ;
			32'h00101adc : data_o = 32'he59256b1 ;
			32'h00101ae0 : data_o = 32'h32781bc0 ;
			32'h00101ae4 : data_o = 32'hf571933e ;
			32'h00101ae8 : data_o = 32'h7817471d ;
			32'h00101aec : data_o = 32'h6658b40c ;
			32'h00101af0 : data_o = 32'hc9998228 ;
			32'h00101af4 : data_o = 32'h59f5ec2b ;
			32'h00101af8 : data_o = 32'hdc008900 ;
			32'h00101afc : data_o = 32'h85481a8c ;
			32'h00101b00 : data_o = 32'h7f7e6981 ;
			32'h00101b04 : data_o = 32'hddcbc828 ;
			32'h00101b08 : data_o = 32'hb2c3c8d6 ;
			32'h00101b0c : data_o = 32'h03a67714 ;
			32'h00101b10 : data_o = 32'h53898d5e ;
			32'h00101b14 : data_o = 32'h1aa16ae3 ;
			32'h00101b18 : data_o = 32'h880fd7e6 ;
			32'h00101b1c : data_o = 32'hc1b6b9c4 ;
			32'h00101b20 : data_o = 32'h16648a19 ;
			32'h00101b24 : data_o = 32'h71e35559 ;
			32'h00101b28 : data_o = 32'h63eaca64 ;
			32'h00101b2c : data_o = 32'h6606d6dc ;
			32'h00101b30 : data_o = 32'h7c08e457 ;
			32'h00101b34 : data_o = 32'h8a572062 ;
			32'h00101b38 : data_o = 32'h7ece0858 ;
			32'h00101b3c : data_o = 32'h26e0878b ;
			32'h00101b40 : data_o = 32'hc37f38a8 ;
			32'h00101b44 : data_o = 32'h0cbbf547 ;
			32'h00101b48 : data_o = 32'hfe24e9ad ;
			32'h00101b4c : data_o = 32'h80d97aad ;
			32'h00101b50 : data_o = 32'h87464a5e ;
			32'h00101b54 : data_o = 32'h5487db47 ;
			32'h00101b58 : data_o = 32'h8622a14d ;
			32'h00101b5c : data_o = 32'h0fd66643 ;
			32'h00101b60 : data_o = 32'h6375f3b4 ;
			32'h00101b64 : data_o = 32'hbdd7e40f ;
			32'h00101b68 : data_o = 32'h59a8e415 ;
			32'h00101b6c : data_o = 32'h78d56c53 ;
			32'h00101b70 : data_o = 32'hd205336f ;
			32'h00101b74 : data_o = 32'hb51e43da ;
			32'h00101b78 : data_o = 32'ha7acbf11 ;
			32'h00101b7c : data_o = 32'h9dc80ab1 ;
			32'h00101b80 : data_o = 32'he510400f ;
			32'h00101b84 : data_o = 32'hf1141d96 ;
			32'h00101b88 : data_o = 32'ha4d8e979 ;
			32'h00101b8c : data_o = 32'h863c497b ;
			32'h00101b90 : data_o = 32'h74733b19 ;
			32'h00101b94 : data_o = 32'h8a349efe ;
			32'h00101b98 : data_o = 32'he693a680 ;
			32'h00101b9c : data_o = 32'hd42b9521 ;
			32'h00101ba0 : data_o = 32'h64a4ef5d ;
			32'h00101ba4 : data_o = 32'h9fb35f88 ;
			32'h00101ba8 : data_o = 32'h6b6b4db8 ;
			32'h00101bac : data_o = 32'hc5cfa1fd ;
			32'h00101bb0 : data_o = 32'h8ed27316 ;
			32'h00101bb4 : data_o = 32'h2e89ed98 ;
			32'h00101bb8 : data_o = 32'he921a5a8 ;
			32'h00101bbc : data_o = 32'hf373e793 ;
			32'h00101bc0 : data_o = 32'hf2a4aaf6 ;
			32'h00101bc4 : data_o = 32'he189d02f ;
			32'h00101bc8 : data_o = 32'h96819705 ;
			32'h00101bcc : data_o = 32'hd11c9032 ;
			32'h00101bd0 : data_o = 32'hff037252 ;
			32'h00101bd4 : data_o = 32'hf97e52dd ;
			32'h00101bd8 : data_o = 32'he0e739a1 ;
			32'h00101bdc : data_o = 32'h8f65295b ;
			32'h00101be0 : data_o = 32'hfc3e747f ;
			32'h00101be4 : data_o = 32'h15c53781 ;
			32'h00101be8 : data_o = 32'h69d1a013 ;
			32'h00101bec : data_o = 32'h84f703a2 ;
			32'h00101bf0 : data_o = 32'hcd3391ec ;
			32'h00101bf4 : data_o = 32'h263a7bbc ;
			32'h00101bf8 : data_o = 32'h3873dbb8 ;
			32'h00101bfc : data_o = 32'hc0f82233 ;
			32'h00101c00 : data_o = 32'h660cf843 ;
			32'h00101c04 : data_o = 32'h5fbd0cf4 ;
			32'h00101c08 : data_o = 32'h3a2299af ;
			32'h00101c0c : data_o = 32'hae26e1a0 ;
			32'h00101c10 : data_o = 32'hb37e3906 ;
			32'h00101c14 : data_o = 32'hae51b5be ;
			32'h00101c18 : data_o = 32'h61e60255 ;
			32'h00101c1c : data_o = 32'h14f51435 ;
			32'h00101c20 : data_o = 32'hae65b1f6 ;
			32'h00101c24 : data_o = 32'h15485b10 ;
			32'h00101c28 : data_o = 32'hf3f503ec ;
			32'h00101c2c : data_o = 32'h9bfd6f6d ;
			32'h00101c30 : data_o = 32'hc6cde1f3 ;
			32'h00101c34 : data_o = 32'hd993f2c0 ;
			32'h00101c38 : data_o = 32'h77cd1c0c ;
			32'h00101c3c : data_o = 32'h7bc64403 ;
			32'h00101c40 : data_o = 32'ha5af03b4 ;
			32'h00101c44 : data_o = 32'h482e6109 ;
			32'h00101c48 : data_o = 32'h413cde96 ;
			32'h00101c4c : data_o = 32'he11a100a ;
			32'h00101c50 : data_o = 32'h73c19225 ;
			32'h00101c54 : data_o = 32'h758e0e0a ;
			32'h00101c58 : data_o = 32'h232bcdb4 ;
			32'h00101c5c : data_o = 32'he72c172c ;
			32'h00101c60 : data_o = 32'h0c3dfe98 ;
			32'h00101c64 : data_o = 32'h35d14d31 ;
			32'h00101c68 : data_o = 32'ha57068be ;
			32'h00101c6c : data_o = 32'ha922533d ;
			32'h00101c70 : data_o = 32'hd0ea9de4 ;
			32'h00101c74 : data_o = 32'ha923561e ;
			32'h00101c78 : data_o = 32'ha8d0d403 ;
			32'h00101c7c : data_o = 32'hbf1664a3 ;
			32'h00101c80 : data_o = 32'hda022658 ;
			32'h00101c84 : data_o = 32'ha42dacb2 ;
			32'h00101c88 : data_o = 32'hc4f62b9b ;
			32'h00101c8c : data_o = 32'hc91951ec ;
			32'h00101c90 : data_o = 32'h1e4e0701 ;
			32'h00101c94 : data_o = 32'h6c6d85f2 ;
			32'h00101c98 : data_o = 32'h76914c75 ;
			32'h00101c9c : data_o = 32'hd7943ae0 ;
			32'h00101ca0 : data_o = 32'ha622dbc5 ;
			32'h00101ca4 : data_o = 32'hdadd5567 ;
			32'h00101ca8 : data_o = 32'h50a2f8ea ;
			32'h00101cac : data_o = 32'h9ab40d44 ;
			32'h00101cb0 : data_o = 32'h43378a9e ;
			32'h00101cb4 : data_o = 32'hd564104f ;
			32'h00101cb8 : data_o = 32'ha9700709 ;
			32'h00101cbc : data_o = 32'h967ad6c5 ;
			32'h00101cc0 : data_o = 32'h18880fda ;
			32'h00101cc4 : data_o = 32'h2d8d0fd8 ;
			32'h00101cc8 : data_o = 32'h1c5bedf5 ;
			32'h00101ccc : data_o = 32'h927a7216 ;
			32'h00101cd0 : data_o = 32'hebda10a6 ;
			32'h00101cd4 : data_o = 32'hb78b0781 ;
			32'h00101cd8 : data_o = 32'h7c682028 ;
			32'h00101cdc : data_o = 32'h4f18f8a1 ;
			32'h00101ce0 : data_o = 32'h296205bb ;
			32'h00101ce4 : data_o = 32'h8ac56baf ;
			32'h00101ce8 : data_o = 32'h98aa9a91 ;
			32'h00101cec : data_o = 32'h654a7297 ;
			32'h00101cf0 : data_o = 32'h410687cb ;
			32'h00101cf4 : data_o = 32'hc8caded1 ;
			32'h00101cf8 : data_o = 32'hc2e9ce67 ;
			32'h00101cfc : data_o = 32'h726ebb4e ;
			32'h00101d00 : data_o = 32'h0583ad00 ;
			32'h00101d04 : data_o = 32'h20d03eac ;
			32'h00101d08 : data_o = 32'haff69a79 ;
			32'h00101d0c : data_o = 32'haf7207dc ;
			32'h00101d10 : data_o = 32'h07c51b01 ;
			32'h00101d14 : data_o = 32'h087f7e4f ;
			32'h00101d18 : data_o = 32'h65d83729 ;
			32'h00101d1c : data_o = 32'hb2e3623e ;
			32'h00101d20 : data_o = 32'hadeba164 ;
			32'h00101d24 : data_o = 32'hc3e56927 ;
			32'h00101d28 : data_o = 32'h96257954 ;
			32'h00101d2c : data_o = 32'hc33ec2ee ;
			32'h00101d30 : data_o = 32'h4e6bb5da ;
			32'h00101d34 : data_o = 32'h37d327ff ;
			32'h00101d38 : data_o = 32'hb8c85291 ;
			32'h00101d3c : data_o = 32'h376440f2 ;
			32'h00101d40 : data_o = 32'hc002b106 ;
			32'h00101d44 : data_o = 32'hc2936b8d ;
			32'h00101d48 : data_o = 32'hcedee57c ;
			32'h00101d4c : data_o = 32'hb992fa64 ;
			32'h00101d50 : data_o = 32'h3144df52 ;
			32'h00101d54 : data_o = 32'hef1a5c9d ;
			32'h00101d58 : data_o = 32'h06f8ece3 ;
			32'h00101d5c : data_o = 32'hb0c0e992 ;
			32'h00101d60 : data_o = 32'hb91a281f ;
			32'h00101d64 : data_o = 32'he6259e52 ;
			32'h00101d68 : data_o = 32'hf28a8ac3 ;
			32'h00101d6c : data_o = 32'he9c873bc ;
			32'h00101d70 : data_o = 32'h0492af6f ;
			32'h00101d74 : data_o = 32'hf23d80aa ;
			32'h00101d78 : data_o = 32'h876826d2 ;
			32'h00101d7c : data_o = 32'h21713904 ;
			32'h00101d80 : data_o = 32'h279f82ca ;
			32'h00101d84 : data_o = 32'h47f7b642 ;
			32'h00101d88 : data_o = 32'h6c509c63 ;
			32'h00101d8c : data_o = 32'h4813c947 ;
			32'h00101d90 : data_o = 32'hb2c303e9 ;
			32'h00101d94 : data_o = 32'h306ca0ea ;
			32'h00101d98 : data_o = 32'h436f3cad ;
			32'h00101d9c : data_o = 32'h424768a1 ;
			32'h00101da0 : data_o = 32'hdde05395 ;
			32'h00101da4 : data_o = 32'h0a8e1c63 ;
			32'h00101da8 : data_o = 32'h79cdf21e ;
			32'h00101dac : data_o = 32'h1e9506cf ;
			32'h00101db0 : data_o = 32'haca0de3e ;
			32'h00101db4 : data_o = 32'h988b1c8f ;
			32'h00101db8 : data_o = 32'he2c10318 ;
			32'h00101dbc : data_o = 32'h4aa1f017 ;
			32'h00101dc0 : data_o = 32'h18036204 ;
			32'h00101dc4 : data_o = 32'h850c10d4 ;
			32'h00101dc8 : data_o = 32'h7fc3fba9 ;
			32'h00101dcc : data_o = 32'h825a1a7e ;
			32'h00101dd0 : data_o = 32'hef63b3a8 ;
			32'h00101dd4 : data_o = 32'hbd5e8491 ;
			32'h00101dd8 : data_o = 32'h1632b2d4 ;
			32'h00101ddc : data_o = 32'h321ca7b5 ;
			32'h00101de0 : data_o = 32'hddc90533 ;
			32'h00101de4 : data_o = 32'h8c2ebef3 ;
			32'h00101de8 : data_o = 32'h6f560757 ;
			32'h00101dec : data_o = 32'h8eb14520 ;
			32'h00101df0 : data_o = 32'hca0514ee ;
			32'h00101df4 : data_o = 32'h6e0b9278 ;
			32'h00101df8 : data_o = 32'hce623e68 ;
			32'h00101dfc : data_o = 32'h3dc2131e ;
			32'h00101e00 : data_o = 32'hd745623a ;
			32'h00101e04 : data_o = 32'h950e811e ;
			32'h00101e08 : data_o = 32'hba65c2e4 ;
			32'h00101e0c : data_o = 32'h1c96a837 ;
			32'h00101e10 : data_o = 32'h0b9310e1 ;
			32'h00101e14 : data_o = 32'h66127f68 ;
			32'h00101e18 : data_o = 32'h75487cd4 ;
			32'h00101e1c : data_o = 32'hfcca073b ;
			32'h00101e20 : data_o = 32'h005c3b45 ;
			32'h00101e24 : data_o = 32'h388b3c9b ;
			32'h00101e28 : data_o = 32'h51bc9ce0 ;
			32'h00101e2c : data_o = 32'hd852f5b2 ;
			32'h00101e30 : data_o = 32'he3882f4e ;
			32'h00101e34 : data_o = 32'hf48aeefd ;
			32'h00101e38 : data_o = 32'h8eb2fbe3 ;
			32'h00101e3c : data_o = 32'h4a2e7284 ;
			32'h00101e40 : data_o = 32'hddada819 ;
			32'h00101e44 : data_o = 32'ha0e61a66 ;
			32'h00101e48 : data_o = 32'hb6f5fda7 ;
			32'h00101e4c : data_o = 32'h40d5524e ;
			32'h00101e50 : data_o = 32'h2a4e7d14 ;
			32'h00101e54 : data_o = 32'h4b7fab84 ;
			32'h00101e58 : data_o = 32'h53766f5d ;
			32'h00101e5c : data_o = 32'hc27e5f5c ;
			32'h00101e60 : data_o = 32'h449afb6b ;
			32'h00101e64 : data_o = 32'hc82400dc ;
			32'h00101e68 : data_o = 32'hfe143fc3 ;
			32'h00101e6c : data_o = 32'hb3176942 ;
			32'h00101e70 : data_o = 32'h703c6742 ;
			32'h00101e74 : data_o = 32'hf2c9da2d ;
			32'h00101e78 : data_o = 32'hac2903c5 ;
			32'h00101e7c : data_o = 32'he49bb6c5 ;
			32'h00101e80 : data_o = 32'hd1a3ec1b ;
			32'h00101e84 : data_o = 32'h8572cc28 ;
			32'h00101e88 : data_o = 32'h41a3e9c1 ;
			32'h00101e8c : data_o = 32'hc595c9f6 ;
			32'h00101e90 : data_o = 32'hdc3212ba ;
			32'h00101e94 : data_o = 32'h30fbe2d9 ;
			32'h00101e98 : data_o = 32'h0c904fd9 ;
			32'h00101e9c : data_o = 32'hfed6b5a8 ;
			32'h00101ea0 : data_o = 32'he152542a ;
			32'h00101ea4 : data_o = 32'h3b40f4f0 ;
			32'h00101ea8 : data_o = 32'h2b3c41f4 ;
			32'h00101eac : data_o = 32'ha7ba82a1 ;
			32'h00101eb0 : data_o = 32'h230d09ae ;
			32'h00101eb4 : data_o = 32'h9389ed37 ;
			32'h00101eb8 : data_o = 32'h2954d134 ;
			32'h00101ebc : data_o = 32'hb83cfaa3 ;
			32'h00101ec0 : data_o = 32'hb32622fc ;
			32'h00101ec4 : data_o = 32'h470fad35 ;
			32'h00101ec8 : data_o = 32'h1f59fcc7 ;
			32'h00101ecc : data_o = 32'hcb7554ec ;
			32'h00101ed0 : data_o = 32'h2fe416e3 ;
			32'h00101ed4 : data_o = 32'hc2b5cf9a ;
			32'h00101ed8 : data_o = 32'he88d2c2b ;
			32'h00101edc : data_o = 32'h101301cd ;
			32'h00101ee0 : data_o = 32'he7f9bb7a ;
			32'h00101ee4 : data_o = 32'hbacc6241 ;
			32'h00101ee8 : data_o = 32'h7e1fa395 ;
			32'h00101eec : data_o = 32'h3e7c621e ;
			32'h00101ef0 : data_o = 32'h148bd859 ;
			32'h00101ef4 : data_o = 32'h74211af6 ;
			32'h00101ef8 : data_o = 32'h5e8a71a8 ;
			32'h00101efc : data_o = 32'hb40afe2c ;
			32'h00101f00 : data_o = 32'hffe1a1ab ;
			32'h00101f04 : data_o = 32'hd019bd6e ;
			32'h00101f08 : data_o = 32'h5ffbeaab ;
			32'h00101f0c : data_o = 32'he7dd3344 ;
			32'h00101f10 : data_o = 32'h235b1f20 ;
			32'h00101f14 : data_o = 32'h9115f0a3 ;
			32'h00101f18 : data_o = 32'h2a9b0398 ;
			32'h00101f1c : data_o = 32'h7639f038 ;
			32'h00101f20 : data_o = 32'h3bce2a56 ;
			32'h00101f24 : data_o = 32'hcf427e3c ;
			32'h00101f28 : data_o = 32'h67a755ee ;
			32'h00101f2c : data_o = 32'h887eadea ;
			32'h00101f30 : data_o = 32'h74e612cd ;
			32'h00101f34 : data_o = 32'hd0c66d1b ;
			32'h00101f38 : data_o = 32'h47f356b4 ;
			32'h00101f3c : data_o = 32'h3662f8dc ;
			32'h00101f40 : data_o = 32'h45469dc5 ;
			32'h00101f44 : data_o = 32'h6037075d ;
			32'h00101f48 : data_o = 32'he9383d62 ;
			32'h00101f4c : data_o = 32'he0caeb3e ;
			32'h00101f50 : data_o = 32'h8ae4f997 ;
			32'h00101f54 : data_o = 32'h19f215d4 ;
			32'h00101f58 : data_o = 32'hbea7c79e ;
			32'h00101f5c : data_o = 32'h77b2cff3 ;
			32'h00101f60 : data_o = 32'h3c424a11 ;
			32'h00101f64 : data_o = 32'h766ee258 ;
			32'h00101f68 : data_o = 32'h0c30b733 ;
			32'h00101f6c : data_o = 32'hd91f2613 ;
			32'h00101f70 : data_o = 32'h4728d5d6 ;
			32'h00101f74 : data_o = 32'h939b9178 ;
			32'h00101f78 : data_o = 32'h8516b929 ;
			32'h00101f7c : data_o = 32'h3d45d583 ;
			32'h00101f80 : data_o = 32'h913a1bb3 ;
			32'h00101f84 : data_o = 32'h8a28afb7 ;
			32'h00101f88 : data_o = 32'h73ae909e ;
			32'h00101f8c : data_o = 32'hda63d15f ;
			32'h00101f90 : data_o = 32'ha996b0f4 ;
			32'h00101f94 : data_o = 32'h74960c98 ;
			32'h00101f98 : data_o = 32'he3c21a43 ;
			32'h00101f9c : data_o = 32'h1f2cd477 ;
			32'h00101fa0 : data_o = 32'h29d7dafe ;
			32'h00101fa4 : data_o = 32'h4791dfca ;
			32'h00101fa8 : data_o = 32'h406ebb11 ;
			32'h00101fac : data_o = 32'hd0091a90 ;
			32'h00101fb0 : data_o = 32'h8d8293db ;
			32'h00101fb4 : data_o = 32'h3cf205a4 ;
			32'h00101fb8 : data_o = 32'h05e55e99 ;
			32'h00101fbc : data_o = 32'hfd617c1b ;
			32'h00101fc0 : data_o = 32'hd1a228c2 ;
			32'h00101fc4 : data_o = 32'h41cfd5f3 ;
			32'h00101fc8 : data_o = 32'h731578d4 ;
			32'h00101fcc : data_o = 32'h93610271 ;
			32'h00101fd0 : data_o = 32'h118fa7e5 ;
			32'h00101fd4 : data_o = 32'h22d11ab7 ;
			32'h00101fd8 : data_o = 32'hdf3d4e3f ;
			32'h00101fdc : data_o = 32'hbf73032a ;
			32'h00101fe0 : data_o = 32'h3425347d ;
			32'h00101fe4 : data_o = 32'h02b21cd1 ;
			32'h00101fe8 : data_o = 32'h79c7e9f3 ;
			32'h00101fec : data_o = 32'h97ad3b67 ;
			32'h00101ff0 : data_o = 32'h49f993cb ;
			32'h00101ff4 : data_o = 32'h01f02566 ;
			32'h00101ff8 : data_o = 32'haacda05b ;
			32'h00101ffc : data_o = 32'habbb3fc1 ;
			32'h00102000 : data_o = 32'ha0bb9932 ;
			32'h00102004 : data_o = 32'h796bd43f ;
			32'h00102008 : data_o = 32'h36b31027 ;
			32'h0010200c : data_o = 32'hbb3f0698 ;
			32'h00102010 : data_o = 32'h5cb761b0 ;
			32'h00102014 : data_o = 32'h9ef69629 ;
			32'h00102018 : data_o = 32'hc73aaae8 ;
			32'h0010201c : data_o = 32'h75b1322e ;
			32'h00102020 : data_o = 32'h2e3af26e ;
			32'h00102024 : data_o = 32'h8e19d5b2 ;
			32'h00102028 : data_o = 32'h02c46522 ;
			32'h0010202c : data_o = 32'hd6351173 ;
			32'h00102030 : data_o = 32'h99009a9f ;
			32'h00102034 : data_o = 32'h7e6b4e2c ;
			32'h00102038 : data_o = 32'h55f50094 ;
			32'h0010203c : data_o = 32'h3f817fca ;
			32'h00102040 : data_o = 32'h3d7f12c6 ;
			32'h00102044 : data_o = 32'hbab9e8ab ;
			32'h00102048 : data_o = 32'h1d1a0cce ;
			32'h0010204c : data_o = 32'hd367bf9e ;
			32'h00102050 : data_o = 32'h2b90fe39 ;
			32'h00102054 : data_o = 32'h00ff6022 ;
			32'h00102058 : data_o = 32'h8d04b718 ;
			32'h0010205c : data_o = 32'hdbd6afa6 ;
			32'h00102060 : data_o = 32'h8905098e ;
			32'h00102064 : data_o = 32'h357e9bd5 ;
			32'h00102068 : data_o = 32'h893718e5 ;
			32'h0010206c : data_o = 32'hf2bffb5b ;
			32'h00102070 : data_o = 32'hc571efe1 ;
			32'h00102074 : data_o = 32'h59030919 ;
			32'h00102078 : data_o = 32'hbf333c84 ;
			32'h0010207c : data_o = 32'h1f50bba3 ;
			32'h00102080 : data_o = 32'hd46a07ad ;
			32'h00102084 : data_o = 32'h5ebdcd85 ;
			32'h00102088 : data_o = 32'h1f54efdb ;
			32'h0010208c : data_o = 32'hdbf8d2a0 ;
			32'h00102090 : data_o = 32'h6129b133 ;
			32'h00102094 : data_o = 32'h86656905 ;
			32'h00102098 : data_o = 32'h41feaff0 ;
			32'h0010209c : data_o = 32'h06bcb11a ;
			32'h001020a0 : data_o = 32'h03628f1d ;
			32'h001020a4 : data_o = 32'hfd62dae5 ;
			32'h001020a8 : data_o = 32'hd22282f4 ;
			32'h001020ac : data_o = 32'ha83ca65e ;
			32'h001020b0 : data_o = 32'h7fa11f0e ;
			32'h001020b4 : data_o = 32'h1291f3bc ;
			32'h001020b8 : data_o = 32'h5048101f ;
			32'h001020bc : data_o = 32'ha891112d ;
			32'h001020c0 : data_o = 32'h5a0e6378 ;
			32'h001020c4 : data_o = 32'h6c22b2a8 ;
			32'h001020c8 : data_o = 32'hcb5cef53 ;
			32'h001020cc : data_o = 32'he701c9ba ;
			32'h001020d0 : data_o = 32'h980551a9 ;
			32'h001020d4 : data_o = 32'h0c33f51b ;
			32'h001020d8 : data_o = 32'hde977a93 ;
			32'h001020dc : data_o = 32'h73ef8672 ;
			32'h001020e0 : data_o = 32'h91cdd408 ;
			32'h001020e4 : data_o = 32'hbae7eb50 ;
			32'h001020e8 : data_o = 32'h937219b5 ;
			32'h001020ec : data_o = 32'h71fe57d9 ;
			32'h001020f0 : data_o = 32'hbea5824b ;
			32'h001020f4 : data_o = 32'h5edddb4d ;
			32'h001020f8 : data_o = 32'hd420df12 ;
			32'h001020fc : data_o = 32'h9ce7f68c ;
			32'h00102100 : data_o = 32'h65b1d08d ;
			32'h00102104 : data_o = 32'h4e9e466c ;
			32'h00102108 : data_o = 32'h4ba91963 ;
			32'h0010210c : data_o = 32'h4a27ebc8 ;
			32'h00102110 : data_o = 32'h8bcae4c3 ;
			32'h00102114 : data_o = 32'h77df899e ;
			32'h00102118 : data_o = 32'h7528787e ;
			32'h0010211c : data_o = 32'h6d90c516 ;
			32'h00102120 : data_o = 32'h6483a39a ;
			32'h00102124 : data_o = 32'hef008580 ;
			32'h00102128 : data_o = 32'h4a28d243 ;
			32'h0010212c : data_o = 32'h632af3c0 ;
			32'h00102130 : data_o = 32'h2815a254 ;
			32'h00102134 : data_o = 32'haadd8c9d ;
			32'h00102138 : data_o = 32'h57ce1561 ;
			32'h0010213c : data_o = 32'h836045aa ;
			32'h00102140 : data_o = 32'h7598c5d1 ;
			32'h00102144 : data_o = 32'h40af8885 ;
			32'h00102148 : data_o = 32'hbeebd801 ;
			32'h0010214c : data_o = 32'h5c3f971c ;
			32'h00102150 : data_o = 32'h330f30a5 ;
			32'h00102154 : data_o = 32'h49f74541 ;
			32'h00102158 : data_o = 32'h096fec60 ;
			32'h0010215c : data_o = 32'he851952e ;
			32'h00102160 : data_o = 32'h3ec6d5e7 ;
			32'h00102164 : data_o = 32'h7332a517 ;
			32'h00102168 : data_o = 32'h530adea9 ;
			32'h0010216c : data_o = 32'hb6000970 ;
			32'h00102170 : data_o = 32'h19feccae ;
			32'h00102174 : data_o = 32'h8a6c03b9 ;
			32'h00102178 : data_o = 32'hefa31d61 ;
			32'h0010217c : data_o = 32'h20b9d9ec ;
			32'h00102180 : data_o = 32'h461f8750 ;
			32'h00102184 : data_o = 32'h4c71ac4a ;
			32'h00102188 : data_o = 32'hfa723ec1 ;
			32'h0010218c : data_o = 32'ha903d838 ;
			32'h00102190 : data_o = 32'hc6213f6a ;
			32'h00102194 : data_o = 32'h0f762e0f ;
			32'h00102198 : data_o = 32'h4e2d948e ;
			32'h0010219c : data_o = 32'hb20d1cc5 ;
			32'h001021a0 : data_o = 32'h2f5f11c1 ;
			32'h001021a4 : data_o = 32'h1d5cca83 ;
			32'h001021a8 : data_o = 32'h8806d605 ;
			32'h001021ac : data_o = 32'h43f79313 ;
			32'h001021b0 : data_o = 32'h9dd2f33e ;
			32'h001021b4 : data_o = 32'h1c15dc5b ;
			32'h001021b8 : data_o = 32'hbb9e6056 ;
			32'h001021bc : data_o = 32'h46731f57 ;
			32'h001021c0 : data_o = 32'hc391f014 ;
			32'h001021c4 : data_o = 32'h67ec7235 ;
			32'h001021c8 : data_o = 32'hd0433831 ;
			32'h001021cc : data_o = 32'hca6ac68a ;
			32'h001021d0 : data_o = 32'ha9810421 ;
			32'h001021d4 : data_o = 32'h6ed1139a ;
			32'h001021d8 : data_o = 32'hb17e877c ;
			32'h001021dc : data_o = 32'hf5c8b187 ;
			32'h001021e0 : data_o = 32'h01a74724 ;
			32'h001021e4 : data_o = 32'h278cd3bb ;
			32'h001021e8 : data_o = 32'h43faf0ba ;
			32'h001021ec : data_o = 32'hdc8bcf25 ;
			32'h001021f0 : data_o = 32'h06bf9326 ;
			32'h001021f4 : data_o = 32'hb83e1ad6 ;
			32'h001021f8 : data_o = 32'h3c4c8c86 ;
			32'h001021fc : data_o = 32'he915124e ;
			32'h00102200 : data_o = 32'hc58687a4 ;
			32'h00102204 : data_o = 32'ha6cae2ef ;
			32'h00102208 : data_o = 32'h5f9f36a9 ;
			32'h0010220c : data_o = 32'h88f4ec85 ;
			32'h00102210 : data_o = 32'h4040aec4 ;
			32'h00102214 : data_o = 32'h15eea129 ;
			32'h00102218 : data_o = 32'h0a93ee8f ;
			32'h0010221c : data_o = 32'h3b78f5d2 ;
			32'h00102220 : data_o = 32'h11924956 ;
			32'h00102224 : data_o = 32'h306960da ;
			32'h00102228 : data_o = 32'hc1e0dba5 ;
			32'h0010222c : data_o = 32'hc8756da6 ;
			32'h00102230 : data_o = 32'h1f3b02f6 ;
			32'h00102234 : data_o = 32'h510e641e ;
			32'h00102238 : data_o = 32'h8cb8dfc2 ;
			32'h0010223c : data_o = 32'hfdd620e9 ;
			32'h00102240 : data_o = 32'he292da6b ;
			32'h00102244 : data_o = 32'he27501e2 ;
			32'h00102248 : data_o = 32'hf5abff38 ;
			32'h0010224c : data_o = 32'h7bcb9a89 ;
			32'h00102250 : data_o = 32'haa5d15b1 ;
			32'h00102254 : data_o = 32'h76777873 ;
			32'h00102258 : data_o = 32'h1d23d645 ;
			32'h0010225c : data_o = 32'h3a5a7854 ;
			32'h00102260 : data_o = 32'hf4a08cf2 ;
			32'h00102264 : data_o = 32'h46bff614 ;
			32'h00102268 : data_o = 32'hc8a7f628 ;
			32'h0010226c : data_o = 32'hb457ab5f ;
			32'h00102270 : data_o = 32'h338c8ef1 ;
			32'h00102274 : data_o = 32'h2bcde46f ;
			32'h00102278 : data_o = 32'hb84b3d3a ;
			32'h0010227c : data_o = 32'h05f7a65d ;
			32'h00102280 : data_o = 32'h9bdcfe0c ;
			32'h00102284 : data_o = 32'hd7e27674 ;
			32'h00102288 : data_o = 32'hd2a945f9 ;
			32'h0010228c : data_o = 32'heaa8f51c ;
			32'h00102290 : data_o = 32'h670c0bd1 ;
			32'h00102294 : data_o = 32'hfe99fcb8 ;
			32'h00102298 : data_o = 32'hea81fdba ;
			32'h0010229c : data_o = 32'h3ac5918b ;
			32'h001022a0 : data_o = 32'hcedc9cef ;
			32'h001022a4 : data_o = 32'he0c2aee5 ;
			32'h001022a8 : data_o = 32'h7b487de2 ;
			32'h001022ac : data_o = 32'hfc783674 ;
			32'h001022b0 : data_o = 32'h12ded76c ;
			32'h001022b4 : data_o = 32'h2d129f4e ;
			32'h001022b8 : data_o = 32'hf76d6753 ;
			32'h001022bc : data_o = 32'had809f90 ;
			32'h001022c0 : data_o = 32'h0cf89208 ;
			32'h001022c4 : data_o = 32'he400d7b4 ;
			32'h001022c8 : data_o = 32'h6d8d5777 ;
			32'h001022cc : data_o = 32'h15de4504 ;
			32'h001022d0 : data_o = 32'hbf6ce736 ;
			32'h001022d4 : data_o = 32'h37a4e23f ;
			32'h001022d8 : data_o = 32'h79a23997 ;
			32'h001022dc : data_o = 32'h065fe098 ;
			32'h001022e0 : data_o = 32'h41942926 ;
			32'h001022e4 : data_o = 32'hfda2056d ;
			32'h001022e8 : data_o = 32'h7f1dba1e ;
			32'h001022ec : data_o = 32'h4308da01 ;
			32'h001022f0 : data_o = 32'heae22c6c ;
			32'h001022f4 : data_o = 32'h5c0d483b ;
			32'h001022f8 : data_o = 32'hd0ea4d03 ;
			32'h001022fc : data_o = 32'hd10d454a ;
			32'h00102300 : data_o = 32'h45fe8ac4 ;
			32'h00102304 : data_o = 32'h100f25ce ;
			32'h00102308 : data_o = 32'ha27d08fd ;
			32'h0010230c : data_o = 32'h791687c1 ;
			32'h00102310 : data_o = 32'hecbc0b77 ;
			32'h00102314 : data_o = 32'h2e0b6279 ;
			32'h00102318 : data_o = 32'h6761754a ;
			32'h0010231c : data_o = 32'hd4064625 ;
			32'h00102320 : data_o = 32'h0f9dc336 ;
			32'h00102324 : data_o = 32'h720eb12d ;
			32'h00102328 : data_o = 32'haf4c4106 ;
			32'h0010232c : data_o = 32'h2bbd2df1 ;
			32'h00102330 : data_o = 32'hac5fb84f ;
			32'h00102334 : data_o = 32'h9854efda ;
			32'h00102338 : data_o = 32'ha2d3054c ;
			32'h0010233c : data_o = 32'h235da150 ;
			32'h00102340 : data_o = 32'hfa979384 ;
			32'h00102344 : data_o = 32'hc573e97e ;
			32'h00102348 : data_o = 32'h01cd4dea ;
			32'h0010234c : data_o = 32'h871e4afd ;
			32'h00102350 : data_o = 32'h0b848e8d ;
			32'h00102354 : data_o = 32'hb435cf8e ;
			32'h00102358 : data_o = 32'h04d6ad32 ;
			32'h0010235c : data_o = 32'h8f0ce71c ;
			32'h00102360 : data_o = 32'hddff093d ;
			32'h00102364 : data_o = 32'h9738b12c ;
			32'h00102368 : data_o = 32'h5915c35a ;
			32'h0010236c : data_o = 32'h7ba5f872 ;
			32'h00102370 : data_o = 32'h971a25f2 ;
			32'h00102374 : data_o = 32'h1982a34d ;
			32'h00102378 : data_o = 32'ha5d89060 ;
			32'h0010237c : data_o = 32'ha73ca2e2 ;
			32'h00102380 : data_o = 32'h74ed574b ;
			32'h00102384 : data_o = 32'h0f01bd24 ;
			32'h00102388 : data_o = 32'h000b00f1 ;
			32'h0010238c : data_o = 32'h0223da8e ;
			32'h00102390 : data_o = 32'h8090b1e0 ;
			32'h00102394 : data_o = 32'h4f4cab60 ;
			32'h00102398 : data_o = 32'hecedf139 ;
			32'h0010239c : data_o = 32'hb9fbb10b ;
			32'h001023a0 : data_o = 32'hb0cb6d4c ;
			32'h001023a4 : data_o = 32'h7e1f59f4 ;
			32'h001023a8 : data_o = 32'h74b62de0 ;
			32'h001023ac : data_o = 32'hc5a495db ;
			32'h001023b0 : data_o = 32'hec1431ff ;
			32'h001023b4 : data_o = 32'h3a527065 ;
			32'h001023b8 : data_o = 32'hbb2c0a67 ;
			32'h001023bc : data_o = 32'ha9c9a882 ;
			32'h001023c0 : data_o = 32'hedfd79a0 ;
			32'h001023c4 : data_o = 32'h710f22a9 ;
			32'h001023c8 : data_o = 32'hf3ca56f0 ;
			32'h001023cc : data_o = 32'hacd85fba ;
			32'h001023d0 : data_o = 32'h1f1407a7 ;
			32'h001023d4 : data_o = 32'h55bb2130 ;
			32'h001023d8 : data_o = 32'hc8d8a899 ;
			32'h001023dc : data_o = 32'h44b79603 ;
			32'h001023e0 : data_o = 32'h0ddaaec8 ;
			32'h001023e4 : data_o = 32'hc146382a ;
			32'h001023e8 : data_o = 32'h0e5a556f ;
			32'h001023ec : data_o = 32'he6fb78eb ;
			32'h001023f0 : data_o = 32'hfe7207c7 ;
			32'h001023f4 : data_o = 32'h37d660f4 ;
			32'h001023f8 : data_o = 32'h8b7ee7df ;
			32'h001023fc : data_o = 32'h711c25cd ;
			32'h00102400 : data_o = 32'ha327c882 ;
			32'h00102404 : data_o = 32'h52c72cc9 ;
			32'h00102408 : data_o = 32'hd37e8c00 ;
			32'h0010240c : data_o = 32'hd7a882a0 ;
			32'h00102410 : data_o = 32'he91af605 ;
			32'h00102414 : data_o = 32'h5b941c04 ;
			32'h00102418 : data_o = 32'h5f84ee0a ;
			32'h0010241c : data_o = 32'h212781d8 ;
			32'h00102420 : data_o = 32'h74d99265 ;
			32'h00102424 : data_o = 32'h1fba0a19 ;
			32'h00102428 : data_o = 32'hcc53c757 ;
			32'h0010242c : data_o = 32'h8cdf6a30 ;
			32'h00102430 : data_o = 32'hf8906a16 ;
			32'h00102434 : data_o = 32'h8dd3f3cd ;
			32'h00102438 : data_o = 32'h6fbc214f ;
			32'h0010243c : data_o = 32'heaea5de2 ;
			32'h00102440 : data_o = 32'h49545f50 ;
			32'h00102444 : data_o = 32'hc7b4e596 ;
			32'h00102448 : data_o = 32'hab323811 ;
			32'h0010244c : data_o = 32'h36fb86e3 ;
			32'h00102450 : data_o = 32'h52be4580 ;
			32'h00102454 : data_o = 32'h261bfb81 ;
			32'h00102458 : data_o = 32'he8066d98 ;
			32'h0010245c : data_o = 32'hbb557191 ;
			32'h00102460 : data_o = 32'h9b3e4b84 ;
			32'h00102464 : data_o = 32'h76889fce ;
			32'h00102468 : data_o = 32'he57e5b67 ;
			32'h0010246c : data_o = 32'hd8b05bbc ;
			32'h00102470 : data_o = 32'hca0d1c01 ;
			32'h00102474 : data_o = 32'h8ecd5b22 ;
			32'h00102478 : data_o = 32'h5936f249 ;
			32'h0010247c : data_o = 32'hf7f31c1b ;
			32'h00102480 : data_o = 32'h6aed94d1 ;
			32'h00102484 : data_o = 32'hfabde366 ;
			32'h00102488 : data_o = 32'h4bde303a ;
			32'h0010248c : data_o = 32'h9a0c2a97 ;
			32'h00102490 : data_o = 32'h66d534f4 ;
			32'h00102494 : data_o = 32'h88ffd269 ;
			32'h00102498 : data_o = 32'hf0dfee90 ;
			32'h0010249c : data_o = 32'hd8535766 ;
			32'h001024a0 : data_o = 32'hf427e1b1 ;
			32'h001024a4 : data_o = 32'h7de8b61d ;
			32'h001024a8 : data_o = 32'h3fa0a615 ;
			32'h001024ac : data_o = 32'hdf009cec ;
			32'h001024b0 : data_o = 32'h9b516520 ;
			32'h001024b4 : data_o = 32'h4f6f1ff8 ;
			32'h001024b8 : data_o = 32'h9a112797 ;
			32'h001024bc : data_o = 32'hda8c15c8 ;
			32'h001024c0 : data_o = 32'h21c12820 ;
			32'h001024c4 : data_o = 32'h1bbc91e6 ;
			32'h001024c8 : data_o = 32'ha54cc162 ;
			32'h001024cc : data_o = 32'h0ee5020c ;
			32'h001024d0 : data_o = 32'h07e02732 ;
			32'h001024d4 : data_o = 32'hd93aa0de ;
			32'h001024d8 : data_o = 32'h9fbec9aa ;
			32'h001024dc : data_o = 32'hde8f057c ;
			32'h001024e0 : data_o = 32'hcb1be91c ;
			32'h001024e4 : data_o = 32'hb5f80229 ;
			32'h001024e8 : data_o = 32'h55d37a84 ;
			32'h001024ec : data_o = 32'h88fd44af ;
			32'h001024f0 : data_o = 32'h3a36602a ;
			32'h001024f4 : data_o = 32'h69dc18f5 ;
			32'h001024f8 : data_o = 32'hcb55c970 ;
			32'h001024fc : data_o = 32'h95d180ed ;
			32'h00102500 : data_o = 32'h997be8e4 ;
			32'h00102504 : data_o = 32'hda7a0537 ;
			32'h00102508 : data_o = 32'h7c09533f ;
			32'h0010250c : data_o = 32'h1952ed3a ;
			32'h00102510 : data_o = 32'hc3e75c43 ;
			32'h00102514 : data_o = 32'h2b3a4149 ;
			32'h00102518 : data_o = 32'h55eba0a4 ;
			32'h0010251c : data_o = 32'h090f102e ;
			32'h00102520 : data_o = 32'h89feeeef ;
			32'h00102524 : data_o = 32'h1cded64d ;
			32'h00102528 : data_o = 32'h735b1d6d ;
			32'h0010252c : data_o = 32'h4ffce502 ;
			32'h00102530 : data_o = 32'h084229a3 ;
			32'h00102534 : data_o = 32'hcd1d42a0 ;
			32'h00102538 : data_o = 32'h0034c1d1 ;
			32'h0010253c : data_o = 32'hbb4bcfa6 ;
			32'h00102540 : data_o = 32'hcbbe9d8c ;
			32'h00102544 : data_o = 32'h35f83ee0 ;
			32'h00102548 : data_o = 32'h23feccc9 ;
			32'h0010254c : data_o = 32'hda15a5dd ;
			32'h00102550 : data_o = 32'hb6623cf2 ;
			32'h00102554 : data_o = 32'h08ec1e6b ;
			32'h00102558 : data_o = 32'hffba3e79 ;
			32'h0010255c : data_o = 32'h52aebb09 ;
			32'h00102560 : data_o = 32'h74fc8ae8 ;
			32'h00102564 : data_o = 32'h5450d7ef ;
			32'h00102568 : data_o = 32'h2b230369 ;
			32'h0010256c : data_o = 32'h6fbbb4c8 ;
			32'h00102570 : data_o = 32'h9063c499 ;
			32'h00102574 : data_o = 32'hcede116e ;
			32'h00102578 : data_o = 32'haf3051d8 ;
			32'h0010257c : data_o = 32'h81cf4ec9 ;
			32'h00102580 : data_o = 32'h03708751 ;
			32'h00102584 : data_o = 32'h43aea268 ;
			32'h00102588 : data_o = 32'h40f53699 ;
			32'h0010258c : data_o = 32'hbbc0417a ;
			32'h00102590 : data_o = 32'hb88efa63 ;
			32'h00102594 : data_o = 32'h4f263050 ;
			32'h00102598 : data_o = 32'ha2007678 ;
			32'h0010259c : data_o = 32'ha11be740 ;
			32'h001025a0 : data_o = 32'h604b41e6 ;
			32'h001025a4 : data_o = 32'h1d278dfc ;
			32'h001025a8 : data_o = 32'h893a204a ;
			32'h001025ac : data_o = 32'hbc2032fb ;
			32'h001025b0 : data_o = 32'hd5284a10 ;
			32'h001025b4 : data_o = 32'hd6be449f ;
			32'h001025b8 : data_o = 32'h952dbf28 ;
			32'h001025bc : data_o = 32'h7ac95411 ;
			32'h001025c0 : data_o = 32'h48cc79db ;
			32'h001025c4 : data_o = 32'h53b91670 ;
			32'h001025c8 : data_o = 32'h3a77f0e3 ;
			32'h001025cc : data_o = 32'h733e5e59 ;
			32'h001025d0 : data_o = 32'h2678de3a ;
			32'h001025d4 : data_o = 32'h5f28c46d ;
			32'h001025d8 : data_o = 32'h5ea7fc0c ;
			32'h001025dc : data_o = 32'h648089c5 ;
			32'h001025e0 : data_o = 32'hffb4fca7 ;
			32'h001025e4 : data_o = 32'h6a6492e4 ;
			32'h001025e8 : data_o = 32'h28fa419e ;
			32'h001025ec : data_o = 32'h6ecf3bb3 ;
			32'h001025f0 : data_o = 32'h91ccfcbc ;
			32'h001025f4 : data_o = 32'hf43b3d5d ;
			32'h001025f8 : data_o = 32'h6f0c2e6c ;
			32'h001025fc : data_o = 32'haaf4c7a6 ;
			32'h00102600 : data_o = 32'ha0f6b0bb ;
			32'h00102604 : data_o = 32'h9fb28ca3 ;
			32'h00102608 : data_o = 32'ha4c9f0d9 ;
			32'h0010260c : data_o = 32'h5d94e8cc ;
			32'h00102610 : data_o = 32'hbbe9fd48 ;
			32'h00102614 : data_o = 32'h1876cd56 ;
			32'h00102618 : data_o = 32'h5248583b ;
			32'h0010261c : data_o = 32'h3651242b ;
			32'h00102620 : data_o = 32'h3348239a ;
			32'h00102624 : data_o = 32'h56814fe3 ;
			32'h00102628 : data_o = 32'h090b4630 ;
			32'h0010262c : data_o = 32'h6096ff4e ;
			32'h00102630 : data_o = 32'h76d755c8 ;
			32'h00102634 : data_o = 32'h03485256 ;
			32'h00102638 : data_o = 32'h31a321d9 ;
			32'h0010263c : data_o = 32'h9981b6bd ;
			32'h00102640 : data_o = 32'he3e092ae ;
			32'h00102644 : data_o = 32'hd78b4039 ;
			32'h00102648 : data_o = 32'h9d776200 ;
			32'h0010264c : data_o = 32'h85d76321 ;
			32'h00102650 : data_o = 32'h81c45a7f ;
			32'h00102654 : data_o = 32'hfca25c91 ;
			32'h00102658 : data_o = 32'hd44c27dc ;
			32'h0010265c : data_o = 32'h287f3378 ;
			32'h00102660 : data_o = 32'h7853b6cd ;
			32'h00102664 : data_o = 32'h69c3e03a ;
			32'h00102668 : data_o = 32'h60793bc2 ;
			32'h0010266c : data_o = 32'hd95f33ee ;
			32'h00102670 : data_o = 32'hcb5f054a ;
			32'h00102674 : data_o = 32'h782dfa1d ;
			32'h00102678 : data_o = 32'h678c390f ;
			32'h0010267c : data_o = 32'h47c1355e ;
			32'h00102680 : data_o = 32'hc538d6a2 ;
			32'h00102684 : data_o = 32'h04a8cefd ;
			32'h00102688 : data_o = 32'h43fd82aa ;
			32'h0010268c : data_o = 32'hc8f578c9 ;
			32'h00102690 : data_o = 32'h2400e2a6 ;
			32'h00102694 : data_o = 32'h37bf7441 ;
			32'h00102698 : data_o = 32'hf427726b ;
			32'h0010269c : data_o = 32'h1adaa64c ;
			32'h001026a0 : data_o = 32'hf81d250d ;
			32'h001026a4 : data_o = 32'hc14373d7 ;
			32'h001026a8 : data_o = 32'haf4b2d28 ;
			32'h001026ac : data_o = 32'hf558a4ed ;
			32'h001026b0 : data_o = 32'hb2e01acf ;
			32'h001026b4 : data_o = 32'hebc0949a ;
			32'h001026b8 : data_o = 32'h058886b0 ;
			32'h001026bc : data_o = 32'h8622f9d2 ;
			32'h001026c0 : data_o = 32'h85520d31 ;
			32'h001026c4 : data_o = 32'hf56183dc ;
			32'h001026c8 : data_o = 32'h0a961d10 ;
			32'h001026cc : data_o = 32'h2c911a04 ;
			32'h001026d0 : data_o = 32'h11ac3192 ;
			32'h001026d4 : data_o = 32'h0a19f45c ;
			32'h001026d8 : data_o = 32'habafca08 ;
			32'h001026dc : data_o = 32'he736a377 ;
			32'h001026e0 : data_o = 32'ha2cf485c ;
			32'h001026e4 : data_o = 32'h0a35200b ;
			32'h001026e8 : data_o = 32'h4ad81968 ;
			32'h001026ec : data_o = 32'h8a0f8eea ;
			32'h001026f0 : data_o = 32'h2aecf781 ;
			32'h001026f4 : data_o = 32'h5526c30c ;
			32'h001026f8 : data_o = 32'h173a92e9 ;
			32'h001026fc : data_o = 32'hf6e0ef6b ;
			32'h00102700 : data_o = 32'hd242648e ;
			32'h00102704 : data_o = 32'h0b52701c ;
			32'h00102708 : data_o = 32'hf40f6cdf ;
			32'h0010270c : data_o = 32'hc2608fe4 ;
			32'h00102710 : data_o = 32'h46ed8902 ;
			32'h00102714 : data_o = 32'h6babd32e ;
			32'h00102718 : data_o = 32'h35b052c4 ;
			32'h0010271c : data_o = 32'h7d0cd25b ;
			32'h00102720 : data_o = 32'h1ff1b834 ;
			32'h00102724 : data_o = 32'h49eb2658 ;
			32'h00102728 : data_o = 32'h217ecf46 ;
			32'h0010272c : data_o = 32'h54f0902b ;
			32'h00102730 : data_o = 32'h1d0ca01c ;
			32'h00102734 : data_o = 32'ha6c4424f ;
			32'h00102738 : data_o = 32'h05e688a1 ;
			32'h0010273c : data_o = 32'he0a7c5b2 ;
			32'h00102740 : data_o = 32'ha3b19805 ;
			32'h00102744 : data_o = 32'h308b0ae3 ;
			32'h00102748 : data_o = 32'hd1fe1dfc ;
			32'h0010274c : data_o = 32'h84da4dea ;
			32'h00102750 : data_o = 32'h2c95b395 ;
			32'h00102754 : data_o = 32'hf3daeede ;
			32'h00102758 : data_o = 32'h582b13d3 ;
			32'h0010275c : data_o = 32'h4325f128 ;
			32'h00102760 : data_o = 32'h6590ddb0 ;
			32'h00102764 : data_o = 32'h165a15e2 ;
			32'h00102768 : data_o = 32'hc82c7006 ;
			32'h0010276c : data_o = 32'h0c50a122 ;
			32'h00102770 : data_o = 32'hc9ff3f98 ;
			32'h00102774 : data_o = 32'h8d3b969f ;
			32'h00102778 : data_o = 32'h9345e7be ;
			32'h0010277c : data_o = 32'h5e225a3f ;
			32'h00102780 : data_o = 32'h7c41e56e ;
			32'h00102784 : data_o = 32'h18aa6e22 ;
			32'h00102788 : data_o = 32'h0542351a ;
			32'h0010278c : data_o = 32'h20c5e3b6 ;
			32'h00102790 : data_o = 32'hf2ed1f70 ;
			32'h00102794 : data_o = 32'h3e970dd7 ;
			32'h00102798 : data_o = 32'h8315d17d ;
			32'h0010279c : data_o = 32'ha5abe6f7 ;
			32'h001027a0 : data_o = 32'h744fb391 ;
			32'h001027a4 : data_o = 32'h19567fb4 ;
			32'h001027a8 : data_o = 32'h29a146e3 ;
			32'h001027ac : data_o = 32'hd0fd488b ;
			32'h001027b0 : data_o = 32'h80746751 ;
			32'h001027b4 : data_o = 32'h1db22124 ;
			32'h001027b8 : data_o = 32'h1427047e ;
			32'h001027bc : data_o = 32'h5ea31eda ;
			32'h001027c0 : data_o = 32'hf4047373 ;
			32'h001027c4 : data_o = 32'hab2cca14 ;
			32'h001027c8 : data_o = 32'h78dfa33a ;
			32'h001027cc : data_o = 32'h5fc8255f ;
			32'h001027d0 : data_o = 32'h6742bdcb ;
			32'h001027d4 : data_o = 32'he1df42d1 ;
			32'h001027d8 : data_o = 32'he416199e ;
			32'h001027dc : data_o = 32'h297a4037 ;
			32'h001027e0 : data_o = 32'h5ac8054d ;
			32'h001027e4 : data_o = 32'h41d14bea ;
			32'h001027e8 : data_o = 32'hc51af548 ;
			32'h001027ec : data_o = 32'hccb869d2 ;
			32'h001027f0 : data_o = 32'h4e99f409 ;
			32'h001027f4 : data_o = 32'h4808daa6 ;
			32'h001027f8 : data_o = 32'h9b09ea60 ;
			32'h001027fc : data_o = 32'hde7da69c ;
			32'h00102800 : data_o = 32'hcb315158 ;
			32'h00102804 : data_o = 32'hdf436702 ;
			32'h00102808 : data_o = 32'ha69f0976 ;
			32'h0010280c : data_o = 32'hc4f6ffce ;
			32'h00102810 : data_o = 32'hb4df5129 ;
			32'h00102814 : data_o = 32'h789cc6d2 ;
			32'h00102818 : data_o = 32'h42b0bd4d ;
			32'h0010281c : data_o = 32'h8cbdea58 ;
			32'h00102820 : data_o = 32'h2bb986ae ;
			32'h00102824 : data_o = 32'h59d0e408 ;
			32'h00102828 : data_o = 32'h5ade7733 ;
			32'h0010282c : data_o = 32'h6b0a72d6 ;
			32'h00102830 : data_o = 32'hd317ffd8 ;
			32'h00102834 : data_o = 32'h2e3f30f2 ;
			32'h00102838 : data_o = 32'he5933276 ;
			32'h0010283c : data_o = 32'h60009e97 ;
			32'h00102840 : data_o = 32'h336f5f1e ;
			32'h00102844 : data_o = 32'h7d8fb761 ;
			32'h00102848 : data_o = 32'hf799b2d2 ;
			32'h0010284c : data_o = 32'h0e6b573b ;
			32'h00102850 : data_o = 32'h88083c0c ;
			32'h00102854 : data_o = 32'heaf4b662 ;
			32'h00102858 : data_o = 32'hbd0979f0 ;
			32'h0010285c : data_o = 32'h7a58cf40 ;
			32'h00102860 : data_o = 32'h4892c640 ;
			32'h00102864 : data_o = 32'h216b8296 ;
			32'h00102868 : data_o = 32'hd4c8c8e2 ;
			32'h0010286c : data_o = 32'h9e3409c0 ;
			32'h00102870 : data_o = 32'hc0335fe1 ;
			32'h00102874 : data_o = 32'he074861e ;
			32'h00102878 : data_o = 32'h64487875 ;
			32'h0010287c : data_o = 32'h81f21aee ;
			32'h00102880 : data_o = 32'hcb4a9ccc ;
			32'h00102884 : data_o = 32'h16a8b294 ;
			32'h00102888 : data_o = 32'h9f3eb675 ;
			32'h0010288c : data_o = 32'h20592d72 ;
			32'h00102890 : data_o = 32'hf3c75669 ;
			32'h00102894 : data_o = 32'h585e7dbc ;
			32'h00102898 : data_o = 32'h0a5e1676 ;
			32'h0010289c : data_o = 32'h92898a97 ;
			32'h001028a0 : data_o = 32'hcf551f96 ;
			32'h001028a4 : data_o = 32'h16a33005 ;
			32'h001028a8 : data_o = 32'h0f53a931 ;
			32'h001028ac : data_o = 32'hce66bd01 ;
			32'h001028b0 : data_o = 32'h2bbf6400 ;
			32'h001028b4 : data_o = 32'hfd2ae019 ;
			32'h001028b8 : data_o = 32'h74226bfb ;
			32'h001028bc : data_o = 32'ha6c01429 ;
			32'h001028c0 : data_o = 32'h3d0ae5ef ;
			32'h001028c4 : data_o = 32'h43fe8058 ;
			32'h001028c8 : data_o = 32'h8ab88bda ;
			32'h001028cc : data_o = 32'h95ebc0ac ;
			32'h001028d0 : data_o = 32'h043db42b ;
			32'h001028d4 : data_o = 32'h8e2d9432 ;
			32'h001028d8 : data_o = 32'h6322ac42 ;
			32'h001028dc : data_o = 32'hb2d01f52 ;
			32'h001028e0 : data_o = 32'hdc611f80 ;
			32'h001028e4 : data_o = 32'hc3ec4a56 ;
			32'h001028e8 : data_o = 32'h9cad8d1a ;
			32'h001028ec : data_o = 32'he3b06a94 ;
			32'h001028f0 : data_o = 32'hc68990cb ;
			32'h001028f4 : data_o = 32'h45ad45ab ;
			32'h001028f8 : data_o = 32'h6e6df7d1 ;
			32'h001028fc : data_o = 32'h72d37032 ;
			32'h00102900 : data_o = 32'h8a036cc0 ;
			32'h00102904 : data_o = 32'hba35740f ;
			32'h00102908 : data_o = 32'hfb301999 ;
			32'h0010290c : data_o = 32'h09e2cb5d ;
			32'h00102910 : data_o = 32'h0ceb38d3 ;
			32'h00102914 : data_o = 32'h57d0ef5f ;
			32'h00102918 : data_o = 32'h90b12191 ;
			32'h0010291c : data_o = 32'h031dd8e1 ;
			32'h00102920 : data_o = 32'hbd022354 ;
			32'h00102924 : data_o = 32'h132fd3d7 ;
			32'h00102928 : data_o = 32'h51c14f45 ;
			32'h0010292c : data_o = 32'h1db958c8 ;
			32'h00102930 : data_o = 32'h80ccd989 ;
			32'h00102934 : data_o = 32'h59ba11b8 ;
			32'h00102938 : data_o = 32'hcbacbc2d ;
			32'h0010293c : data_o = 32'h73aef6d6 ;
			32'h00102940 : data_o = 32'h20a4077f ;
			32'h00102944 : data_o = 32'hb9871b86 ;
			32'h00102948 : data_o = 32'h9eda3f42 ;
			32'h0010294c : data_o = 32'h11d26dc5 ;
			32'h00102950 : data_o = 32'h9934726b ;
			32'h00102954 : data_o = 32'h985b6216 ;
			32'h00102958 : data_o = 32'h12099206 ;
			32'h0010295c : data_o = 32'hd53667f0 ;
			32'h00102960 : data_o = 32'h174ad049 ;
			32'h00102964 : data_o = 32'h500ec1fb ;
			32'h00102968 : data_o = 32'he60e0e17 ;
			32'h0010296c : data_o = 32'hb5c858b0 ;
			32'h00102970 : data_o = 32'h97b3886b ;
			32'h00102974 : data_o = 32'h1324c0a8 ;
			32'h00102978 : data_o = 32'h5e717cd1 ;
			32'h0010297c : data_o = 32'h662f28c2 ;
			32'h00102980 : data_o = 32'h55bf15c6 ;
			32'h00102984 : data_o = 32'hd1806b2e ;
			32'h00102988 : data_o = 32'h9d9b7b68 ;
			32'h0010298c : data_o = 32'hd3b41c6d ;
			32'h00102990 : data_o = 32'hcbd9af5e ;
			32'h00102994 : data_o = 32'h710f9735 ;
			32'h00102998 : data_o = 32'hd7b288bc ;
			32'h0010299c : data_o = 32'h07b2fc81 ;
			32'h001029a0 : data_o = 32'h9a4c161d ;
			32'h001029a4 : data_o = 32'h161283b9 ;
			32'h001029a8 : data_o = 32'h9e7bc388 ;
			32'h001029ac : data_o = 32'h977dfb8a ;
			32'h001029b0 : data_o = 32'he1a5a510 ;
			32'h001029b4 : data_o = 32'h08e5f282 ;
			32'h001029b8 : data_o = 32'h807d197c ;
			32'h001029bc : data_o = 32'h133bfa2d ;
			32'h001029c0 : data_o = 32'h1b4cf683 ;
			32'h001029c4 : data_o = 32'h1a449ecd ;
			32'h001029c8 : data_o = 32'h3298d6a9 ;
			32'h001029cc : data_o = 32'h420f7869 ;
			32'h001029d0 : data_o = 32'hae9e3af8 ;
			32'h001029d4 : data_o = 32'h8686b739 ;
			32'h001029d8 : data_o = 32'he11c4081 ;
			32'h001029dc : data_o = 32'h9bf18e65 ;
			32'h001029e0 : data_o = 32'h098ec46d ;
			32'h001029e4 : data_o = 32'h5af80746 ;
			32'h001029e8 : data_o = 32'h9f6d60d6 ;
			32'h001029ec : data_o = 32'h0e52fd24 ;
			32'h001029f0 : data_o = 32'h30a001ea ;
			32'h001029f4 : data_o = 32'hb9041aec ;
			32'h001029f8 : data_o = 32'hf7c050c7 ;
			32'h001029fc : data_o = 32'h4654ecd8 ;
			32'h00102a00 : data_o = 32'h01ec3a4d ;
			32'h00102a04 : data_o = 32'hb56c3663 ;
			32'h00102a08 : data_o = 32'h36553714 ;
			32'h00102a0c : data_o = 32'h3aa1f35a ;
			32'h00102a10 : data_o = 32'h68b444fd ;
			32'h00102a14 : data_o = 32'hcb9f7bc8 ;
			32'h00102a18 : data_o = 32'h7c95a431 ;
			32'h00102a1c : data_o = 32'h14288832 ;
			32'h00102a20 : data_o = 32'hd3cf8358 ;
			32'h00102a24 : data_o = 32'h57c8753d ;
			32'h00102a28 : data_o = 32'h66bc55c8 ;
			32'h00102a2c : data_o = 32'h486f6489 ;
			32'h00102a30 : data_o = 32'hc039e096 ;
			32'h00102a34 : data_o = 32'h4e14fc1e ;
			32'h00102a38 : data_o = 32'h64e588c7 ;
			32'h00102a3c : data_o = 32'h0a21dc6a ;
			32'h00102a40 : data_o = 32'h53a2bfba ;
			32'h00102a44 : data_o = 32'h4a6bacd6 ;
			32'h00102a48 : data_o = 32'h1a2c9ce9 ;
			32'h00102a4c : data_o = 32'h027efa87 ;
			32'h00102a50 : data_o = 32'h6d1d4d8f ;
			32'h00102a54 : data_o = 32'h242663d9 ;
			32'h00102a58 : data_o = 32'h02782893 ;
			32'h00102a5c : data_o = 32'ha9776566 ;
			32'h00102a60 : data_o = 32'h50b33b9e ;
			32'h00102a64 : data_o = 32'hdb63001e ;
			32'h00102a68 : data_o = 32'h4fd7a407 ;
			32'h00102a6c : data_o = 32'hf78837da ;
			32'h00102a70 : data_o = 32'ha8f5eed9 ;
			32'h00102a74 : data_o = 32'hac21dc78 ;
			32'h00102a78 : data_o = 32'hd1a22592 ;
			32'h00102a7c : data_o = 32'heb505339 ;
			32'h00102a80 : data_o = 32'h84fea8c8 ;
			32'h00102a84 : data_o = 32'h77211004 ;
			32'h00102a88 : data_o = 32'h3498c9e7 ;
			32'h00102a8c : data_o = 32'h57ab64d2 ;
			32'h00102a90 : data_o = 32'hb7224e1b ;
			32'h00102a94 : data_o = 32'h47287ed4 ;
			32'h00102a98 : data_o = 32'h9c40ed02 ;
			32'h00102a9c : data_o = 32'hd56ee243 ;
			32'h00102aa0 : data_o = 32'h884120d2 ;
			32'h00102aa4 : data_o = 32'h028518b3 ;
			32'h00102aa8 : data_o = 32'h5836b52a ;
			32'h00102aac : data_o = 32'heaef4114 ;
			32'h00102ab0 : data_o = 32'h2048eb24 ;
			32'h00102ab4 : data_o = 32'h6403b04a ;
			32'h00102ab8 : data_o = 32'he382c611 ;
			32'h00102abc : data_o = 32'h03064cb6 ;
			32'h00102ac0 : data_o = 32'h384c054e ;
			32'h00102ac4 : data_o = 32'h9a341909 ;
			32'h00102ac8 : data_o = 32'h3ff54f9d ;
			32'h00102acc : data_o = 32'h2df36729 ;
			32'h00102ad0 : data_o = 32'h3ab15bd3 ;
			32'h00102ad4 : data_o = 32'h3ad65060 ;
			32'h00102ad8 : data_o = 32'h3426cb53 ;
			32'h00102adc : data_o = 32'h8ff8ffe9 ;
			32'h00102ae0 : data_o = 32'h003f93dc ;
			32'h00102ae4 : data_o = 32'h09c81756 ;
			32'h00102ae8 : data_o = 32'hff780d21 ;
			32'h00102aec : data_o = 32'hb9480b80 ;
			32'h00102af0 : data_o = 32'h4d0ded28 ;
			32'h00102af4 : data_o = 32'h90072497 ;
			32'h00102af8 : data_o = 32'h1843a442 ;
			32'h00102afc : data_o = 32'h5b9eb4f7 ;
			32'h00102b00 : data_o = 32'h8724fd6c ;
			32'h00102b04 : data_o = 32'h6f044235 ;
			32'h00102b08 : data_o = 32'h1da82e27 ;
			32'h00102b0c : data_o = 32'h21c99aff ;
			32'h00102b10 : data_o = 32'hab7917e6 ;
			32'h00102b14 : data_o = 32'h8523f92f ;
			32'h00102b18 : data_o = 32'h6d4980c7 ;
			32'h00102b1c : data_o = 32'h5678f92a ;
			32'h00102b20 : data_o = 32'hf153a39a ;
			32'h00102b24 : data_o = 32'hd215312e ;
			32'h00102b28 : data_o = 32'he5a2bf4e ;
			32'h00102b2c : data_o = 32'h63c6d3bf ;
			32'h00102b30 : data_o = 32'h905118c6 ;
			32'h00102b34 : data_o = 32'h96cfc405 ;
			32'h00102b38 : data_o = 32'h2d2cbc55 ;
			32'h00102b3c : data_o = 32'h9138eb2f ;
			32'h00102b40 : data_o = 32'h3c6d158d ;
			32'h00102b44 : data_o = 32'h32a58303 ;
			32'h00102b48 : data_o = 32'h9237463d ;
			32'h00102b4c : data_o = 32'hfc8dd8b8 ;
			32'h00102b50 : data_o = 32'hde6b3ff1 ;
			32'h00102b54 : data_o = 32'h8309ccce ;
			32'h00102b58 : data_o = 32'h88467be1 ;
			32'h00102b5c : data_o = 32'h63ab5909 ;
			32'h00102b60 : data_o = 32'h8fd4e319 ;
			32'h00102b64 : data_o = 32'hf1bc1d13 ;
			32'h00102b68 : data_o = 32'h44e3c60a ;
			32'h00102b6c : data_o = 32'h94ca15d3 ;
			32'h00102b70 : data_o = 32'h7a5f80be ;
			32'h00102b74 : data_o = 32'h2ef9ed45 ;
			32'h00102b78 : data_o = 32'h5a45a00a ;
			32'h00102b7c : data_o = 32'h7fc39c0e ;
			32'h00102b80 : data_o = 32'h2be9ad67 ;
			32'h00102b84 : data_o = 32'h266fe9e2 ;
			32'h00102b88 : data_o = 32'h8e4c1086 ;
			32'h00102b8c : data_o = 32'hf210e31f ;
			32'h00102b90 : data_o = 32'h5f34c134 ;
			32'h00102b94 : data_o = 32'h071217cb ;
			32'h00102b98 : data_o = 32'h401f98e9 ;
			32'h00102b9c : data_o = 32'h9527efc2 ;
			32'h00102ba0 : data_o = 32'h355d18ee ;
			32'h00102ba4 : data_o = 32'hd1e5e08b ;
			32'h00102ba8 : data_o = 32'h09d1d64d ;
			32'h00102bac : data_o = 32'hb3e43e47 ;
			32'h00102bb0 : data_o = 32'hecb36a50 ;
			32'h00102bb4 : data_o = 32'h6b24be2a ;
			32'h00102bb8 : data_o = 32'hf6f11e65 ;
			32'h00102bbc : data_o = 32'ha1ac389e ;
			32'h00102bc0 : data_o = 32'h1252bac6 ;
			32'h00102bc4 : data_o = 32'hcfbc6f30 ;
			32'h00102bc8 : data_o = 32'hd19240c1 ;
			32'h00102bcc : data_o = 32'h0a0e6b54 ;
			32'h00102bd0 : data_o = 32'h15c52b77 ;
			32'h00102bd4 : data_o = 32'hc5769881 ;
			32'h00102bd8 : data_o = 32'h1e930ee6 ;
			32'h00102bdc : data_o = 32'hb8ca4fbe ;
			32'h00102be0 : data_o = 32'heb1d5355 ;
			32'h00102be4 : data_o = 32'h263527a8 ;
			32'h00102be8 : data_o = 32'hc13250d1 ;
			32'h00102bec : data_o = 32'hf53ca836 ;
			32'h00102bf0 : data_o = 32'h611d33b1 ;
			32'h00102bf4 : data_o = 32'h3e2ac359 ;
			32'h00102bf8 : data_o = 32'hfb7fd69e ;
			32'h00102bfc : data_o = 32'h74e89351 ;
			32'h00102c00 : data_o = 32'h361a0040 ;
			32'h00102c04 : data_o = 32'h1f897e8b ;
			32'h00102c08 : data_o = 32'h572cb91d ;
			32'h00102c0c : data_o = 32'he35112da ;
			32'h00102c10 : data_o = 32'h2b4f30e8 ;
			32'h00102c14 : data_o = 32'h52fb12fb ;
			32'h00102c18 : data_o = 32'hfae7f5fb ;
			32'h00102c1c : data_o = 32'hd83a7efa ;
			32'h00102c20 : data_o = 32'hf4afad3c ;
			32'h00102c24 : data_o = 32'hcee55c4b ;
			32'h00102c28 : data_o = 32'h00ae66b0 ;
			32'h00102c2c : data_o = 32'h6090db78 ;
			32'h00102c30 : data_o = 32'h892d3f9d ;
			32'h00102c34 : data_o = 32'h2c3d120e ;
			32'h00102c38 : data_o = 32'h6095367e ;
			32'h00102c3c : data_o = 32'hcc888851 ;
			32'h00102c40 : data_o = 32'h7a01b0e3 ;
			32'h00102c44 : data_o = 32'hd71e4b1d ;
			32'h00102c48 : data_o = 32'hc0e6acde ;
			32'h00102c4c : data_o = 32'h152f2d0e ;
			32'h00102c50 : data_o = 32'hb9d16622 ;
			32'h00102c54 : data_o = 32'he1532d8c ;
			32'h00102c58 : data_o = 32'h82fcfa2f ;
			32'h00102c5c : data_o = 32'h22eee580 ;
			32'h00102c60 : data_o = 32'h81fb5a5f ;
			32'h00102c64 : data_o = 32'h51ecf0b6 ;
			32'h00102c68 : data_o = 32'h4325b208 ;
			32'h00102c6c : data_o = 32'h235b0ec1 ;
			32'h00102c70 : data_o = 32'h3329a088 ;
			32'h00102c74 : data_o = 32'h1a09bb79 ;
			32'h00102c78 : data_o = 32'h6e79fb7c ;
			32'h00102c7c : data_o = 32'h6ed26ab2 ;
			32'h00102c80 : data_o = 32'h82fc33e5 ;
			32'h00102c84 : data_o = 32'h1879570a ;
			32'h00102c88 : data_o = 32'h2d0d436c ;
			32'h00102c8c : data_o = 32'h90e70d76 ;
			32'h00102c90 : data_o = 32'h1ddbeb2a ;
			32'h00102c94 : data_o = 32'h1d42f0e3 ;
			32'h00102c98 : data_o = 32'hd128e20a ;
			32'h00102c9c : data_o = 32'h16b1cf25 ;
			32'h00102ca0 : data_o = 32'h58993c80 ;
			32'h00102ca4 : data_o = 32'h3f8eeeb3 ;
			32'h00102ca8 : data_o = 32'h0df8d2af ;
			32'h00102cac : data_o = 32'h8b34ffbf ;
			32'h00102cb0 : data_o = 32'hbf875c10 ;
			32'h00102cb4 : data_o = 32'h1866c4a9 ;
			32'h00102cb8 : data_o = 32'h9ca42066 ;
			32'h00102cbc : data_o = 32'hce090410 ;
			32'h00102cc0 : data_o = 32'heba15f0c ;
			32'h00102cc4 : data_o = 32'h7d800d6d ;
			32'h00102cc8 : data_o = 32'hcd053e84 ;
			32'h00102ccc : data_o = 32'h1d99636e ;
			32'h00102cd0 : data_o = 32'h33b7c2bc ;
			32'h00102cd4 : data_o = 32'haa79efc4 ;
			32'h00102cd8 : data_o = 32'hb65b88ff ;
			32'h00102cdc : data_o = 32'h144c2b6e ;
			32'h00102ce0 : data_o = 32'hda24f9e0 ;
			32'h00102ce4 : data_o = 32'hfb8fa4ca ;
			32'h00102ce8 : data_o = 32'h20c834a4 ;
			32'h00102cec : data_o = 32'hf75ebde2 ;
			32'h00102cf0 : data_o = 32'h848e19d7 ;
			32'h00102cf4 : data_o = 32'h4f331d19 ;
			32'h00102cf8 : data_o = 32'h21e65c26 ;
			32'h00102cfc : data_o = 32'h30f4dc4c ;
			32'h00102d00 : data_o = 32'h39ed0dc4 ;
			32'h00102d04 : data_o = 32'hc17a2ec4 ;
			32'h00102d08 : data_o = 32'h76d1c537 ;
			32'h00102d0c : data_o = 32'h7f5b7eeb ;
			32'h00102d10 : data_o = 32'h56753b20 ;
			32'h00102d14 : data_o = 32'h923d9d84 ;
			32'h00102d18 : data_o = 32'hc363c9a4 ;
			32'h00102d1c : data_o = 32'h0ee5736f ;
			32'h00102d20 : data_o = 32'h203670c2 ;
			32'h00102d24 : data_o = 32'h04c9aa75 ;
			32'h00102d28 : data_o = 32'h1f423c7c ;
			32'h00102d2c : data_o = 32'hec978c58 ;
			32'h00102d30 : data_o = 32'h9b1ba3a5 ;
			32'h00102d34 : data_o = 32'hbd2dc9e7 ;
			32'h00102d38 : data_o = 32'h5ac7bd6b ;
			32'h00102d3c : data_o = 32'h6d9fa5df ;
			32'h00102d40 : data_o = 32'habf6ce01 ;
			32'h00102d44 : data_o = 32'h1618ab96 ;
			32'h00102d48 : data_o = 32'h65ae4989 ;
			32'h00102d4c : data_o = 32'h0dde4b99 ;
			32'h00102d50 : data_o = 32'hb9a061fe ;
			32'h00102d54 : data_o = 32'h9efcf1e1 ;
			32'h00102d58 : data_o = 32'h6db8c66e ;
			32'h00102d5c : data_o = 32'h77a9751c ;
			32'h00102d60 : data_o = 32'h3b030630 ;
			32'h00102d64 : data_o = 32'h68985f1c ;
			32'h00102d68 : data_o = 32'haa673575 ;
			32'h00102d6c : data_o = 32'h30e8131d ;
			32'h00102d70 : data_o = 32'h9dbaea4d ;
			32'h00102d74 : data_o = 32'h90472503 ;
			32'h00102d78 : data_o = 32'hed1fa3fa ;
			32'h00102d7c : data_o = 32'hf5217b45 ;
			32'h00102d80 : data_o = 32'hed0fdc63 ;
			32'h00102d84 : data_o = 32'h2afd9c7b ;
			32'h00102d88 : data_o = 32'he9c31112 ;
			32'h00102d8c : data_o = 32'hec491289 ;
			32'h00102d90 : data_o = 32'h6db9c4c7 ;
			32'h00102d94 : data_o = 32'ha7f96584 ;
			32'h00102d98 : data_o = 32'h5375955c ;
			32'h00102d9c : data_o = 32'hbaf2c12c ;
			32'h00102da0 : data_o = 32'h9fd64fe3 ;
			32'h00102da4 : data_o = 32'h86e8b49f ;
			32'h00102da8 : data_o = 32'hee044ddc ;
			32'h00102dac : data_o = 32'h671c2d6d ;
			32'h00102db0 : data_o = 32'h000d7e3e ;
			32'h00102db4 : data_o = 32'h0ce514fd ;
			32'h00102db8 : data_o = 32'h78d3f906 ;
			32'h00102dbc : data_o = 32'hb4df1b00 ;
			32'h00102dc0 : data_o = 32'h021d5c5b ;
			32'h00102dc4 : data_o = 32'hd74e38f4 ;
			32'h00102dc8 : data_o = 32'h7e1fb96f ;
			32'h00102dcc : data_o = 32'hdacf7fc3 ;
			32'h00102dd0 : data_o = 32'h5a2c1fee ;
			32'h00102dd4 : data_o = 32'h1647a3eb ;
			32'h00102dd8 : data_o = 32'h60a6fe31 ;
			32'h00102ddc : data_o = 32'h83402984 ;
			32'h00102de0 : data_o = 32'h85753ce1 ;
			32'h00102de4 : data_o = 32'h2bd2c3c3 ;
			32'h00102de8 : data_o = 32'h093a7250 ;
			32'h00102dec : data_o = 32'ha0c60477 ;
			32'h00102df0 : data_o = 32'h96f6ef81 ;
			32'h00102df4 : data_o = 32'h7010e3b0 ;
			32'h00102df8 : data_o = 32'h0e2bcc2d ;
			32'h00102dfc : data_o = 32'h57d4a44c ;
			32'h00102e00 : data_o = 32'h37d4baef ;
			32'h00102e04 : data_o = 32'h14dd19fe ;
			32'h00102e08 : data_o = 32'ha54f83e4 ;
			32'h00102e0c : data_o = 32'hdd127510 ;
			32'h00102e10 : data_o = 32'h6f27dae1 ;
			32'h00102e14 : data_o = 32'h5601fc93 ;
			32'h00102e18 : data_o = 32'h0b860003 ;
			32'h00102e1c : data_o = 32'hbea454d6 ;
			32'h00102e20 : data_o = 32'h1afec75d ;
			32'h00102e24 : data_o = 32'h500d97f7 ;
			32'h00102e28 : data_o = 32'hefee1f3a ;
			32'h00102e2c : data_o = 32'h8dc31dc5 ;
			32'h00102e30 : data_o = 32'h9aa6494d ;
			32'h00102e34 : data_o = 32'h9e55467e ;
			32'h00102e38 : data_o = 32'h76405f93 ;
			32'h00102e3c : data_o = 32'h943e549f ;
			32'h00102e40 : data_o = 32'ha23ef578 ;
			32'h00102e44 : data_o = 32'hd22777fc ;
			32'h00102e48 : data_o = 32'he1de8224 ;
			32'h00102e4c : data_o = 32'ha03d4612 ;
			32'h00102e50 : data_o = 32'hd3e664fa ;
			32'h00102e54 : data_o = 32'hd5a06868 ;
			32'h00102e58 : data_o = 32'h4b4444b9 ;
			32'h00102e5c : data_o = 32'h8b7ade0e ;
			32'h00102e60 : data_o = 32'h6e152558 ;
			32'h00102e64 : data_o = 32'h1df70c64 ;
			32'h00102e68 : data_o = 32'hf1d31e6d ;
			32'h00102e6c : data_o = 32'hb508877c ;
			32'h00102e70 : data_o = 32'h1314a881 ;
			32'h00102e74 : data_o = 32'hb20d169e ;
			32'h00102e78 : data_o = 32'hf15a42ef ;
			32'h00102e7c : data_o = 32'h202d81d7 ;
			32'h00102e80 : data_o = 32'hff40280a ;
			32'h00102e84 : data_o = 32'h2fc77e2a ;
			32'h00102e88 : data_o = 32'he9973d9e ;
			32'h00102e8c : data_o = 32'hf6295de4 ;
			32'h00102e90 : data_o = 32'hfa3b03af ;
			32'h00102e94 : data_o = 32'h61742521 ;
			32'h00102e98 : data_o = 32'hddbafa57 ;
			32'h00102e9c : data_o = 32'he26d2d72 ;
			32'h00102ea0 : data_o = 32'he1989180 ;
			32'h00102ea4 : data_o = 32'h9c6abe70 ;
			32'h00102ea8 : data_o = 32'h006a6c89 ;
			32'h00102eac : data_o = 32'h07888520 ;
			32'h00102eb0 : data_o = 32'h8541f0f2 ;
			32'h00102eb4 : data_o = 32'h6d38f30f ;
			32'h00102eb8 : data_o = 32'h4c323d21 ;
			32'h00102ebc : data_o = 32'h064e2712 ;
			32'h00102ec0 : data_o = 32'hed5df7ba ;
			32'h00102ec4 : data_o = 32'h28cb42d4 ;
			32'h00102ec8 : data_o = 32'h63a6a365 ;
			32'h00102ecc : data_o = 32'h3c873cb3 ;
			32'h00102ed0 : data_o = 32'h598ab1d9 ;
			32'h00102ed4 : data_o = 32'h770017a7 ;
			32'h00102ed8 : data_o = 32'h95ffa726 ;
			32'h00102edc : data_o = 32'h9bea3b44 ;
			32'h00102ee0 : data_o = 32'ha1c34e46 ;
			32'h00102ee4 : data_o = 32'h687c89c9 ;
			32'h00102ee8 : data_o = 32'h61b8591f ;
			32'h00102eec : data_o = 32'ha0a1ba5c ;
			32'h00102ef0 : data_o = 32'h886c9865 ;
			32'h00102ef4 : data_o = 32'hf5a18cb6 ;
			32'h00102ef8 : data_o = 32'h01458185 ;
			32'h00102efc : data_o = 32'hca7792af ;
			32'h00102f00 : data_o = 32'h1ab3418c ;
			32'h00102f04 : data_o = 32'h1e9d8740 ;
			32'h00102f08 : data_o = 32'h2d205bc6 ;
			32'h00102f0c : data_o = 32'he929716e ;
			32'h00102f10 : data_o = 32'h7dcc3ab7 ;
			32'h00102f14 : data_o = 32'h91e50f21 ;
			32'h00102f18 : data_o = 32'h406e3f00 ;
			32'h00102f1c : data_o = 32'h7c32f88f ;
			32'h00102f20 : data_o = 32'he23a7546 ;
			32'h00102f24 : data_o = 32'hd532b1d1 ;
			32'h00102f28 : data_o = 32'hcfb1654e ;
			32'h00102f2c : data_o = 32'h58c84901 ;
			32'h00102f30 : data_o = 32'h5523faeb ;
			32'h00102f34 : data_o = 32'h7047903f ;
			32'h00102f38 : data_o = 32'h8f18bece ;
			32'h00102f3c : data_o = 32'hc7d2794a ;
			32'h00102f40 : data_o = 32'h80c489a6 ;
			32'h00102f44 : data_o = 32'h14f2266e ;
			32'h00102f48 : data_o = 32'hfdcbce0f ;
			32'h00102f4c : data_o = 32'h89ae05c9 ;
			32'h00102f50 : data_o = 32'h8f0ec3d0 ;
			32'h00102f54 : data_o = 32'hd2f5e599 ;
			32'h00102f58 : data_o = 32'h89840366 ;
			32'h00102f5c : data_o = 32'hf6b68e5d ;
			32'h00102f60 : data_o = 32'h868990f0 ;
			32'h00102f64 : data_o = 32'h1fc35e47 ;
			32'h00102f68 : data_o = 32'hb3c2a0a3 ;
			32'h00102f6c : data_o = 32'h0a26a117 ;
			32'h00102f70 : data_o = 32'h4c2414c1 ;
			32'h00102f74 : data_o = 32'h2e8bad87 ;
			32'h00102f78 : data_o = 32'h3abc4c7e ;
			32'h00102f7c : data_o = 32'h45f3e537 ;
			32'h00102f80 : data_o = 32'haa2aab36 ;
			32'h00102f84 : data_o = 32'h8dcdf9ae ;
			32'h00102f88 : data_o = 32'h2ebd83c2 ;
			32'h00102f8c : data_o = 32'h8fa5407d ;
			32'h00102f90 : data_o = 32'h0c6e75f3 ;
			32'h00102f94 : data_o = 32'h3e5ab968 ;
			32'h00102f98 : data_o = 32'h6fd74757 ;
			32'h00102f9c : data_o = 32'h2ae1d14a ;
			32'h00102fa0 : data_o = 32'hd6fa0f88 ;
			32'h00102fa4 : data_o = 32'h86c4db68 ;
			32'h00102fa8 : data_o = 32'h6ca6ff75 ;
			32'h00102fac : data_o = 32'h95d0568d ;
			32'h00102fb0 : data_o = 32'h66f4b32c ;
			32'h00102fb4 : data_o = 32'hd333099b ;
			32'h00102fb8 : data_o = 32'hb7b8a77e ;
			32'h00102fbc : data_o = 32'h7cc5f347 ;
			32'h00102fc0 : data_o = 32'ha1bb2108 ;
			32'h00102fc4 : data_o = 32'h88860285 ;
			32'h00102fc8 : data_o = 32'h84c84d06 ;
			32'h00102fcc : data_o = 32'h8fa8a304 ;
			32'h00102fd0 : data_o = 32'hcd54975f ;
			32'h00102fd4 : data_o = 32'h3df67496 ;
			32'h00102fd8 : data_o = 32'hc29a9ac2 ;
			32'h00102fdc : data_o = 32'h862bfc5d ;
			32'h00102fe0 : data_o = 32'h78d7026c ;
			32'h00102fe4 : data_o = 32'h7efdaa58 ;
			32'h00102fe8 : data_o = 32'ha3e894fd ;
			32'h00102fec : data_o = 32'h158b102f ;
			32'h00102ff0 : data_o = 32'hcf3bd67c ;
			32'h00102ff4 : data_o = 32'h106c16f4 ;
			32'h00102ff8 : data_o = 32'h36601363 ;
			32'h00102ffc : data_o = 32'h7b4c159e ;
			32'h00103000 : data_o = 32'h65839bcc ;
			32'h00103004 : data_o = 32'ha66de535 ;
			32'h00103008 : data_o = 32'h030cfb9f ;
			32'h0010300c : data_o = 32'hc0c6496e ;
			32'h00103010 : data_o = 32'h845f63be ;
			32'h00103014 : data_o = 32'h67c17da9 ;
			32'h00103018 : data_o = 32'h583a739d ;
			32'h0010301c : data_o = 32'hcc20f921 ;
			32'h00103020 : data_o = 32'h36691ee9 ;
			32'h00103024 : data_o = 32'h62cf83c7 ;
			32'h00103028 : data_o = 32'hf669be85 ;
			32'h0010302c : data_o = 32'h1c1b764a ;
			32'h00103030 : data_o = 32'he54b6b83 ;
			32'h00103034 : data_o = 32'hf82b86f7 ;
			32'h00103038 : data_o = 32'h60703110 ;
			32'h0010303c : data_o = 32'h61892929 ;
			32'h00103040 : data_o = 32'hb74a9f11 ;
			32'h00103044 : data_o = 32'h3dc0f586 ;
			32'h00103048 : data_o = 32'hd34bb5d5 ;
			32'h0010304c : data_o = 32'hf4198324 ;
			32'h00103050 : data_o = 32'h53388b7f ;
			32'h00103054 : data_o = 32'h1f5c94ed ;
			32'h00103058 : data_o = 32'h3aac0c36 ;
			32'h0010305c : data_o = 32'h8f02d4de ;
			32'h00103060 : data_o = 32'h2f93ac17 ;
			32'h00103064 : data_o = 32'hb526d35b ;
			32'h00103068 : data_o = 32'h5d9b7a4b ;
			32'h0010306c : data_o = 32'hffe95d57 ;
			32'h00103070 : data_o = 32'hf8c79e95 ;
			32'h00103074 : data_o = 32'h212a49f9 ;
			32'h00103078 : data_o = 32'h09f4adb9 ;
			32'h0010307c : data_o = 32'h29fe8113 ;
			32'h00103080 : data_o = 32'ha379d142 ;
			32'h00103084 : data_o = 32'ha95b06bd ;
			32'h00103088 : data_o = 32'h45435845 ;
			32'h0010308c : data_o = 32'h4f495450 ;
			32'h00103090 : data_o = 32'h2121214e ;
			32'h00103094 : data_o = 32'h0000000a ;
			32'h00103098 : data_o = 32'h3d3d3d3d ;
			32'h0010309c : data_o = 32'h3d3d3d3d ;
			32'h001030a0 : data_o = 32'h3d3d3d3d ;
			32'h001030a4 : data_o = 32'h0000000a ;
			32'h001030a8 : data_o = 32'h4350454d ;
			32'h001030ac : data_o = 32'h2020203a ;
			32'h001030b0 : data_o = 32'h00007830 ;
			32'h001030b4 : data_o = 32'h41434d0a ;
			32'h001030b8 : data_o = 32'h3a455355 ;
			32'h001030bc : data_o = 32'h00783020 ;
			32'h001030c0 : data_o = 32'h56544d0a ;
			32'h001030c4 : data_o = 32'h203a4c41 ;
			32'h001030c8 : data_o = 32'h00783020 ;
			32'h001030cc : data_o = 32'h00100000 ;
			default : data_o = 32'h00000000 ;
		endcase 
	end
endmodule
