module rom_1p #(
	int Depth, 
 	int DATA_WIDTH = 32, 
 	int ADDR_WIDTH = 32 
 ) (
	input logic clk_i, 
	input logic req_i, 
	input logic [ADDR_WIDTH-1:0] addr_i, 
	output logic [DATA_WIDTH-1:0] data_o 
 );
	always_ff @(posedge clk_i) begin
		case (addr_i)
			32'h00100000 : data_o = 32'h3c20106f ;
			32'h00100004 : data_o = 32'h3be0106f ;
			32'h00100008 : data_o = 32'h3ba0106f ;
			32'h0010000c : data_o = 32'h3b60106f ;
			32'h00100010 : data_o = 32'h3b20106f ;
			32'h00100014 : data_o = 32'h3ae0106f ;
			32'h00100018 : data_o = 32'h3aa0106f ;
			32'h0010001c : data_o = 32'h3a60106f ;
			32'h00100020 : data_o = 32'h3a20106f ;
			32'h00100024 : data_o = 32'h39e0106f ;
			32'h00100028 : data_o = 32'h39a0106f ;
			32'h0010002c : data_o = 32'h3960106f ;
			32'h00100030 : data_o = 32'h3920106f ;
			32'h00100034 : data_o = 32'h38e0106f ;
			32'h00100038 : data_o = 32'h38a0106f ;
			32'h0010003c : data_o = 32'h3860106f ;
			32'h00100040 : data_o = 32'h3820106f ;
			32'h00100044 : data_o = 32'h0400006f ;
			32'h00100048 : data_o = 32'h37a0106f ;
			32'h0010004c : data_o = 32'h3760106f ;
			32'h00100050 : data_o = 32'h3720106f ;
			32'h00100054 : data_o = 32'h36e0106f ;
			32'h00100058 : data_o = 32'h36a0106f ;
			32'h0010005c : data_o = 32'h3660106f ;
			32'h00100060 : data_o = 32'h3620106f ;
			32'h00100064 : data_o = 32'h35e0106f ;
			32'h00100068 : data_o = 32'h35a0106f ;
			32'h0010006c : data_o = 32'h3560106f ;
			32'h00100070 : data_o = 32'h3520106f ;
			32'h00100074 : data_o = 32'h34e0106f ;
			32'h00100078 : data_o = 32'h34a0106f ;
			32'h0010007c : data_o = 32'h3460106f ;
			32'h00100080 : data_o = 32'h14f0106f ;
			32'h00100084 : data_o = 32'hc686715d ;
			32'h00100088 : data_o = 32'hc29ac496 ;
			32'h0010008c : data_o = 32'hde22c09e ;
			32'h00100090 : data_o = 32'hda2edc2a ;
			32'h00100094 : data_o = 32'hd636d832 ;
			32'h00100098 : data_o = 32'hd23ed43a ;
			32'h0010009c : data_o = 32'hce46d042 ;
			32'h001000a0 : data_o = 32'hca76cc72 ;
			32'h001000a4 : data_o = 32'hc67ec87a ;
			32'h001000a8 : data_o = 32'h10ef0880 ;
			32'h001000ac : data_o = 32'h872a7740 ;
			32'h001000b0 : data_o = 32'h00100797 ;
			32'h001000b4 : data_o = 32'hf5878793 ;
			32'h001000b8 : data_o = 32'h0797c398 ;
			32'h001000bc : data_o = 32'h87930010 ;
			32'h001000c0 : data_o = 32'h4705f527 ;
			32'h001000c4 : data_o = 32'h0001c398 ;
			32'h001000c8 : data_o = 32'h42a640b6 ;
			32'h001000cc : data_o = 32'h43864316 ;
			32'h001000d0 : data_o = 32'h55625472 ;
			32'h001000d4 : data_o = 32'h564255d2 ;
			32'h001000d8 : data_o = 32'h572256b2 ;
			32'h001000dc : data_o = 32'h58025792 ;
			32'h001000e0 : data_o = 32'h4e6248f2 ;
			32'h001000e4 : data_o = 32'h4f424ed2 ;
			32'h001000e8 : data_o = 32'h61614fb2 ;
			32'h001000ec : data_o = 32'h30200073 ;
			32'h001000f0 : data_o = 32'hd6067179 ;
			32'h001000f4 : data_o = 32'h1800d422 ;
			32'h001000f8 : data_o = 32'hfca42e23 ;
			32'h001000fc : data_o = 32'hfe042623 ;
			32'h00100100 : data_o = 32'h2783a005 ;
			32'h00100104 : data_o = 32'h2703fec4 ;
			32'h00100108 : data_o = 32'h97bafdc4 ;
			32'h0010010c : data_o = 32'h0007c783 ;
			32'h00100110 : data_o = 32'h00ef853e ;
			32'h00100114 : data_o = 32'h27837ff0 ;
			32'h00100118 : data_o = 32'h0785fec4 ;
			32'h0010011c : data_o = 32'hfef42623 ;
			32'h00100120 : data_o = 32'hfec42783 ;
			32'h00100124 : data_o = 32'hfdc42703 ;
			32'h00100128 : data_o = 32'hc78397ba ;
			32'h0010012c : data_o = 32'hfbf10007 ;
			32'h00100130 : data_o = 32'h00010001 ;
			32'h00100134 : data_o = 32'h542250b2 ;
			32'h00100138 : data_o = 32'h80826145 ;
			32'h0010013c : data_o = 32'hd6067179 ;
			32'h00100140 : data_o = 32'h1800d422 ;
			32'h00100144 : data_o = 32'hfca42e23 ;
			32'h00100148 : data_o = 32'hfe042623 ;
			32'h0010014c : data_o = 32'h00efa0a1 ;
			32'h00100150 : data_o = 32'h86aa7fd0 ;
			32'h00100154 : data_o = 32'hfec42783 ;
			32'h00100158 : data_o = 32'hfdc42703 ;
			32'h0010015c : data_o = 32'hf71397ba ;
			32'h00100160 : data_o = 32'h80230ff6 ;
			32'h00100164 : data_o = 32'h278300e7 ;
			32'h00100168 : data_o = 32'h2703fec4 ;
			32'h0010016c : data_o = 32'h97bafdc4 ;
			32'h00100170 : data_o = 32'h0007c703 ;
			32'h00100174 : data_o = 32'h1a6347a9 ;
			32'h00100178 : data_o = 32'h278300f7 ;
			32'h0010017c : data_o = 32'h2703fec4 ;
			32'h00100180 : data_o = 32'h97bafdc4 ;
			32'h00100184 : data_o = 32'h00078023 ;
			32'h00100188 : data_o = 32'h2783a005 ;
			32'h0010018c : data_o = 32'h0785fec4 ;
			32'h00100190 : data_o = 32'hfef42623 ;
			32'h00100194 : data_o = 32'hfec42703 ;
			32'h00100198 : data_o = 32'hdae347fd ;
			32'h0010019c : data_o = 32'h2783fae7 ;
			32'h001001a0 : data_o = 32'h07fdfdc4 ;
			32'h001001a4 : data_o = 32'h00078023 ;
			32'h001001a8 : data_o = 32'h542250b2 ;
			32'h001001ac : data_o = 32'h80826145 ;
			32'h001001b0 : data_o = 32'hd6227179 ;
			32'h001001b4 : data_o = 32'h2e231800 ;
			32'h001001b8 : data_o = 32'h2703fca4 ;
			32'h001001bc : data_o = 32'h0793fdc4 ;
			32'h001001c0 : data_o = 32'h07b30640 ;
			32'h001001c4 : data_o = 32'h222302f7 ;
			32'h001001c8 : data_o = 32'h2423fef4 ;
			32'h001001cc : data_o = 32'h2623fe04 ;
			32'h001001d0 : data_o = 32'ha819fe04 ;
			32'h001001d4 : data_o = 32'hfe842783 ;
			32'h001001d8 : data_o = 32'h24230785 ;
			32'h001001dc : data_o = 32'h2783fef4 ;
			32'h001001e0 : data_o = 32'h0785fec4 ;
			32'h001001e4 : data_o = 32'hfef42623 ;
			32'h001001e8 : data_o = 32'hfec42703 ;
			32'h001001ec : data_o = 32'hfe442783 ;
			32'h001001f0 : data_o = 32'hfef762e3 ;
			32'h001001f4 : data_o = 32'hfe842783 ;
			32'h001001f8 : data_o = 32'h5432853e ;
			32'h001001fc : data_o = 32'h80826145 ;
			32'h00100200 : data_o = 32'hd6227179 ;
			32'h00100204 : data_o = 32'h2e231800 ;
			32'h00100208 : data_o = 32'h2c23fca4 ;
			32'h0010020c : data_o = 32'h2a23fcb4 ;
			32'h00100210 : data_o = 32'h2623fcc4 ;
			32'h00100214 : data_o = 32'h2423fe04 ;
			32'h00100218 : data_o = 32'ha8f1fe04 ;
			32'h0010021c : data_o = 32'hfe842783 ;
			32'h00100220 : data_o = 32'h2703078e ;
			32'h00100224 : data_o = 32'h57b3fdc4 ;
			32'h00100228 : data_o = 32'h02a300f7 ;
			32'h0010022c : data_o = 32'h2783fef4 ;
			32'h00100230 : data_o = 32'h078efe84 ;
			32'h00100234 : data_o = 32'hfd442703 ;
			32'h00100238 : data_o = 32'h00074703 ;
			32'h0010023c : data_o = 32'h873e97ba ;
			32'h00100240 : data_o = 32'hfd842783 ;
			32'h00100244 : data_o = 32'hc78397ba ;
			32'h00100248 : data_o = 32'h86be0007 ;
			32'h0010024c : data_o = 32'hfe842783 ;
			32'h00100250 : data_o = 32'h078e0791 ;
			32'h00100254 : data_o = 32'hfd442703 ;
			32'h00100258 : data_o = 32'h47030705 ;
			32'h0010025c : data_o = 32'h97ba0007 ;
			32'h00100260 : data_o = 32'h2783873e ;
			32'h00100264 : data_o = 32'h97bafd84 ;
			32'h00100268 : data_o = 32'h0007c783 ;
			32'h0010026c : data_o = 32'h07c297b6 ;
			32'h00100270 : data_o = 32'h270383c1 ;
			32'h00100274 : data_o = 32'h0721fe84 ;
			32'h00100278 : data_o = 32'h2683070e ;
			32'h0010027c : data_o = 32'h0689fd44 ;
			32'h00100280 : data_o = 32'h0006c683 ;
			32'h00100284 : data_o = 32'h86ba9736 ;
			32'h00100288 : data_o = 32'hfd842703 ;
			32'h0010028c : data_o = 32'h47039736 ;
			32'h00100290 : data_o = 32'h97ba0007 ;
			32'h00100294 : data_o = 32'h83c107c2 ;
			32'h00100298 : data_o = 32'hfe842703 ;
			32'h0010029c : data_o = 32'h070e0731 ;
			32'h001002a0 : data_o = 32'hfd442683 ;
			32'h001002a4 : data_o = 32'hc683068d ;
			32'h001002a8 : data_o = 32'h97360006 ;
			32'h001002ac : data_o = 32'h270386ba ;
			32'h001002b0 : data_o = 32'h9736fd84 ;
			32'h001002b4 : data_o = 32'h00074703 ;
			32'h001002b8 : data_o = 32'h132397ba ;
			32'h001002bc : data_o = 32'h5703fef4 ;
			32'h001002c0 : data_o = 32'h0793fe64 ;
			32'h001002c4 : data_o = 32'hf6630fe0 ;
			32'h001002c8 : data_o = 32'h079300e7 ;
			32'h001002cc : data_o = 32'h13230ff0 ;
			32'h001002d0 : data_o = 32'h4783fef4 ;
			32'h001002d4 : data_o = 32'h07c2fe54 ;
			32'h001002d8 : data_o = 32'h570383c1 ;
			32'h001002dc : data_o = 32'h0763fe64 ;
			32'h001002e0 : data_o = 32'h278300f7 ;
			32'h001002e4 : data_o = 32'h0785fec4 ;
			32'h001002e8 : data_o = 32'hfef42623 ;
			32'h001002ec : data_o = 32'hfe842783 ;
			32'h001002f0 : data_o = 32'h24230785 ;
			32'h001002f4 : data_o = 32'h2703fef4 ;
			32'h001002f8 : data_o = 32'h478dfe84 ;
			32'h001002fc : data_o = 32'hf2e7d0e3 ;
			32'h00100300 : data_o = 32'hfec42783 ;
			32'h00100304 : data_o = 32'h5432853e ;
			32'h00100308 : data_o = 32'h80826145 ;
			32'h0010030c : data_o = 32'hd6227179 ;
			32'h00100310 : data_o = 32'h2e231800 ;
			32'h00100314 : data_o = 32'h2c23fca4 ;
			32'h00100318 : data_o = 32'h2a23fcb4 ;
			32'h0010031c : data_o = 32'h2623fcc4 ;
			32'h00100320 : data_o = 32'h2423fe04 ;
			32'h00100324 : data_o = 32'haa11fe04 ;
			32'h00100328 : data_o = 32'hfe842783 ;
			32'h0010032c : data_o = 32'h2703078e ;
			32'h00100330 : data_o = 32'h57b3fdc4 ;
			32'h00100334 : data_o = 32'h02a300f7 ;
			32'h00100338 : data_o = 32'h2783fef4 ;
			32'h0010033c : data_o = 32'h078efe84 ;
			32'h00100340 : data_o = 32'hfd442703 ;
			32'h00100344 : data_o = 32'h00074703 ;
			32'h00100348 : data_o = 32'h873e97ba ;
			32'h0010034c : data_o = 32'hfd842783 ;
			32'h00100350 : data_o = 32'hc78397ba ;
			32'h00100354 : data_o = 32'h86be0007 ;
			32'h00100358 : data_o = 32'hfe842783 ;
			32'h0010035c : data_o = 32'h078e0791 ;
			32'h00100360 : data_o = 32'hfd442703 ;
			32'h00100364 : data_o = 32'h47030705 ;
			32'h00100368 : data_o = 32'h97ba0007 ;
			32'h0010036c : data_o = 32'h2783873e ;
			32'h00100370 : data_o = 32'h97bafd84 ;
			32'h00100374 : data_o = 32'h0007c783 ;
			32'h00100378 : data_o = 32'h07c297b6 ;
			32'h0010037c : data_o = 32'h270383c1 ;
			32'h00100380 : data_o = 32'h0721fe84 ;
			32'h00100384 : data_o = 32'h2683070e ;
			32'h00100388 : data_o = 32'h0689fd44 ;
			32'h0010038c : data_o = 32'h0006c683 ;
			32'h00100390 : data_o = 32'h86ba9736 ;
			32'h00100394 : data_o = 32'hfd842703 ;
			32'h00100398 : data_o = 32'h47039736 ;
			32'h0010039c : data_o = 32'h97ba0007 ;
			32'h001003a0 : data_o = 32'h83c107c2 ;
			32'h001003a4 : data_o = 32'hfe842703 ;
			32'h001003a8 : data_o = 32'h070e0731 ;
			32'h001003ac : data_o = 32'hfd442683 ;
			32'h001003b0 : data_o = 32'hc683068d ;
			32'h001003b4 : data_o = 32'h97360006 ;
			32'h001003b8 : data_o = 32'h270386ba ;
			32'h001003bc : data_o = 32'h9736fd84 ;
			32'h001003c0 : data_o = 32'h00074703 ;
			32'h001003c4 : data_o = 32'h132397ba ;
			32'h001003c8 : data_o = 32'h5703fef4 ;
			32'h001003cc : data_o = 32'h0793fe64 ;
			32'h001003d0 : data_o = 32'hf6630fe0 ;
			32'h001003d4 : data_o = 32'h079300e7 ;
			32'h001003d8 : data_o = 32'h13230ff0 ;
			32'h001003dc : data_o = 32'h4783fef4 ;
			32'h001003e0 : data_o = 32'h07c2fe54 ;
			32'h001003e4 : data_o = 32'h570383c1 ;
			32'h001003e8 : data_o = 32'h0363fe64 ;
			32'h001003ec : data_o = 32'h478304f7 ;
			32'h001003f0 : data_o = 32'h07c2fe54 ;
			32'h001003f4 : data_o = 32'h570383c1 ;
			32'h001003f8 : data_o = 32'h7f63fe64 ;
			32'h001003fc : data_o = 32'h470300f7 ;
			32'h00100400 : data_o = 32'h5783fe54 ;
			32'h00100404 : data_o = 32'h07b3fe64 ;
			32'h00100408 : data_o = 32'h873e40f7 ;
			32'h0010040c : data_o = 32'hfec42783 ;
			32'h00100410 : data_o = 32'h262397ba ;
			32'h00100414 : data_o = 32'ha829fef4 ;
			32'h00100418 : data_o = 32'hfe645703 ;
			32'h0010041c : data_o = 32'hfe544783 ;
			32'h00100420 : data_o = 32'h40f707b3 ;
			32'h00100424 : data_o = 32'h2783873e ;
			32'h00100428 : data_o = 32'h97bafec4 ;
			32'h0010042c : data_o = 32'hfef42623 ;
			32'h00100430 : data_o = 32'hfe842783 ;
			32'h00100434 : data_o = 32'h24230785 ;
			32'h00100438 : data_o = 32'h2703fef4 ;
			32'h0010043c : data_o = 32'h478dfe84 ;
			32'h00100440 : data_o = 32'heee7d4e3 ;
			32'h00100444 : data_o = 32'hfec42783 ;
			32'h00100448 : data_o = 32'h5432853e ;
			32'h0010044c : data_o = 32'h80826145 ;
			32'h00100450 : data_o = 32'hd6067179 ;
			32'h00100454 : data_o = 32'h1800d422 ;
			32'h00100458 : data_o = 32'hfca42e23 ;
			32'h0010045c : data_o = 32'hfe042623 ;
			32'h00100460 : data_o = 32'h471da8a9 ;
			32'h00100464 : data_o = 32'hfec42783 ;
			32'h00100468 : data_o = 32'h40f707b3 ;
			32'h0010046c : data_o = 32'h2703078a ;
			32'h00100470 : data_o = 32'h57b3fdc4 ;
			32'h00100474 : data_o = 32'hf79300f7 ;
			32'h00100478 : data_o = 32'h8bbd0ff7 ;
			32'h0010047c : data_o = 32'hfef405a3 ;
			32'h00100480 : data_o = 32'hfeb44703 ;
			32'h00100484 : data_o = 32'hec6347a5 ;
			32'h00100488 : data_o = 32'h478300e7 ;
			32'h0010048c : data_o = 32'h8793feb4 ;
			32'h00100490 : data_o = 32'hf7930307 ;
			32'h00100494 : data_o = 32'h853e0ff7 ;
			32'h00100498 : data_o = 32'h479000ef ;
			32'h0010049c : data_o = 32'h4783a811 ;
			32'h001004a0 : data_o = 32'h8793feb4 ;
			32'h001004a4 : data_o = 32'hf7930377 ;
			32'h001004a8 : data_o = 32'h853e0ff7 ;
			32'h001004ac : data_o = 32'h465000ef ;
			32'h001004b0 : data_o = 32'hfec42783 ;
			32'h001004b4 : data_o = 32'h26230785 ;
			32'h001004b8 : data_o = 32'h2703fef4 ;
			32'h001004bc : data_o = 32'h479dfec4 ;
			32'h001004c0 : data_o = 32'hfae7d1e3 ;
			32'h001004c4 : data_o = 32'h00ef4529 ;
			32'h001004c8 : data_o = 32'h000144b0 ;
			32'h001004cc : data_o = 32'h542250b2 ;
			32'h001004d0 : data_o = 32'h80826145 ;
			32'h001004d4 : data_o = 32'hd6067179 ;
			32'h001004d8 : data_o = 32'h1800d422 ;
			32'h001004dc : data_o = 32'hfca42e23 ;
			32'h001004e0 : data_o = 32'hfdc42783 ;
			32'h001004e4 : data_o = 32'hfef42423 ;
			32'h001004e8 : data_o = 32'hfe042623 ;
			32'h001004ec : data_o = 32'h2703a835 ;
			32'h001004f0 : data_o = 32'h47a9fe84 ;
			32'h001004f4 : data_o = 32'h02f777b3 ;
			32'h001004f8 : data_o = 32'h0ff7f793 ;
			32'h001004fc : data_o = 32'h03078793 ;
			32'h00100500 : data_o = 32'h0ff7f713 ;
			32'h00100504 : data_o = 32'hfec42783 ;
			32'h00100508 : data_o = 32'h97a217c1 ;
			32'h0010050c : data_o = 32'hfee78a23 ;
			32'h00100510 : data_o = 32'hfe842703 ;
			32'h00100514 : data_o = 32'h57b347a9 ;
			32'h00100518 : data_o = 32'h242302f7 ;
			32'h0010051c : data_o = 32'h2783fef4 ;
			32'h00100520 : data_o = 32'h0785fec4 ;
			32'h00100524 : data_o = 32'hfef42623 ;
			32'h00100528 : data_o = 32'hfec42703 ;
			32'h0010052c : data_o = 32'hd0e3478d ;
			32'h00100530 : data_o = 32'h478dfce7 ;
			32'h00100534 : data_o = 32'hfef42623 ;
			32'h00100538 : data_o = 32'h2783a839 ;
			32'h0010053c : data_o = 32'h17c1fec4 ;
			32'h00100540 : data_o = 32'hc78397a2 ;
			32'h00100544 : data_o = 32'h853eff47 ;
			32'h00100548 : data_o = 32'h3c9000ef ;
			32'h0010054c : data_o = 32'hfec42783 ;
			32'h00100550 : data_o = 32'h262317fd ;
			32'h00100554 : data_o = 32'h2783fef4 ;
			32'h00100558 : data_o = 32'hd0e3fec4 ;
			32'h0010055c : data_o = 32'h0001fe07 ;
			32'h00100560 : data_o = 32'h50b20001 ;
			32'h00100564 : data_o = 32'h61455422 ;
			32'h00100568 : data_o = 32'h71058082 ;
			32'h0010056c : data_o = 32'h1c112e23 ;
			32'h00100570 : data_o = 32'h1c812c23 ;
			32'h00100574 : data_o = 32'h07b71380 ;
			32'h00100578 : data_o = 32'h47058000 ;
			32'h0010057c : data_o = 32'h1717c398 ;
			32'h00100580 : data_o = 32'h07130000 ;
			32'h00100584 : data_o = 32'h07936de7 ;
			32'h00100588 : data_o = 32'h86baf344 ;
			32'h0010058c : data_o = 32'h08000713 ;
			32'h00100590 : data_o = 32'h85b6863a ;
			32'h00100594 : data_o = 32'h10ef853e ;
			32'h00100598 : data_o = 32'h26234b80 ;
			32'h0010059c : data_o = 32'ha035fe04 ;
			32'h001005a0 : data_o = 32'hfec42783 ;
			32'h001005a4 : data_o = 32'h97a217c1 ;
			32'h001005a8 : data_o = 32'hf447c783 ;
			32'h001005ac : data_o = 32'h03f7f793 ;
			32'h001005b0 : data_o = 32'h0ff7f713 ;
			32'h001005b4 : data_o = 32'hfec42783 ;
			32'h001005b8 : data_o = 32'h97a217c1 ;
			32'h001005bc : data_o = 32'hece78223 ;
			32'h001005c0 : data_o = 32'hfec42783 ;
			32'h001005c4 : data_o = 32'h26230785 ;
			32'h001005c8 : data_o = 32'h2703fef4 ;
			32'h001005cc : data_o = 32'h0793fec4 ;
			32'h001005d0 : data_o = 32'hf7e307f0 ;
			32'h001005d4 : data_o = 32'h2823fce7 ;
			32'h001005d8 : data_o = 32'h57fdea04 ;
			32'h001005dc : data_o = 32'heaf42623 ;
			32'h001005e0 : data_o = 32'hfe0405a3 ;
			32'h001005e4 : data_o = 32'h0523aa2d ;
			32'h001005e8 : data_o = 32'ha205fe04 ;
			32'h001005ec : data_o = 32'hfeb44783 ;
			32'h001005f0 : data_o = 32'hf7938385 ;
			32'h001005f4 : data_o = 32'h97130ff7 ;
			32'h001005f8 : data_o = 32'h47830027 ;
			32'h001005fc : data_o = 32'h97bafea4 ;
			32'h00100600 : data_o = 32'h00179713 ;
			32'h00100604 : data_o = 32'hfeb44783 ;
			32'h00100608 : data_o = 32'h97ba8b85 ;
			32'h0010060c : data_o = 32'h00279713 ;
			32'h00100610 : data_o = 32'hfeb44683 ;
			32'h00100614 : data_o = 32'hfea44783 ;
			32'h00100618 : data_o = 32'h97b6078e ;
			32'h0010061c : data_o = 32'h1741078a ;
			32'h00100620 : data_o = 32'h47039722 ;
			32'h00100624 : data_o = 32'h17c1ec47 ;
			32'h00100628 : data_o = 32'h8e2397a2 ;
			32'h0010062c : data_o = 32'h4783e2e7 ;
			32'h00100630 : data_o = 32'h8385feb4 ;
			32'h00100634 : data_o = 32'h0ff7f793 ;
			32'h00100638 : data_o = 32'h00279713 ;
			32'h0010063c : data_o = 32'hfea44783 ;
			32'h00100640 : data_o = 32'h971397ba ;
			32'h00100644 : data_o = 32'h47830017 ;
			32'h00100648 : data_o = 32'h8b85feb4 ;
			32'h0010064c : data_o = 32'h078a97ba ;
			32'h00100650 : data_o = 32'h00178713 ;
			32'h00100654 : data_o = 32'hfeb44683 ;
			32'h00100658 : data_o = 32'hfea44783 ;
			32'h0010065c : data_o = 32'h97b6078e ;
			32'h00100660 : data_o = 32'h0785078a ;
			32'h00100664 : data_o = 32'h97221741 ;
			32'h00100668 : data_o = 32'hec474703 ;
			32'h0010066c : data_o = 32'h97a217c1 ;
			32'h00100670 : data_o = 32'he2e78e23 ;
			32'h00100674 : data_o = 32'hfeb44783 ;
			32'h00100678 : data_o = 32'hf7938385 ;
			32'h0010067c : data_o = 32'h97130ff7 ;
			32'h00100680 : data_o = 32'h47830027 ;
			32'h00100684 : data_o = 32'h97bafea4 ;
			32'h00100688 : data_o = 32'h00179713 ;
			32'h0010068c : data_o = 32'hfeb44783 ;
			32'h00100690 : data_o = 32'h97ba8b85 ;
			32'h00100694 : data_o = 32'h8713078a ;
			32'h00100698 : data_o = 32'h46830027 ;
			32'h0010069c : data_o = 32'h4783feb4 ;
			32'h001006a0 : data_o = 32'h078efea4 ;
			32'h001006a4 : data_o = 32'h078a97b6 ;
			32'h001006a8 : data_o = 32'h17410789 ;
			32'h001006ac : data_o = 32'h47039722 ;
			32'h001006b0 : data_o = 32'h17c1ec47 ;
			32'h001006b4 : data_o = 32'h8e2397a2 ;
			32'h001006b8 : data_o = 32'h4783e2e7 ;
			32'h001006bc : data_o = 32'h8385feb4 ;
			32'h001006c0 : data_o = 32'h0ff7f793 ;
			32'h001006c4 : data_o = 32'h00279713 ;
			32'h001006c8 : data_o = 32'hfea44783 ;
			32'h001006cc : data_o = 32'h971397ba ;
			32'h001006d0 : data_o = 32'h47830017 ;
			32'h001006d4 : data_o = 32'h8b85feb4 ;
			32'h001006d8 : data_o = 32'h078a97ba ;
			32'h001006dc : data_o = 32'h00378713 ;
			32'h001006e0 : data_o = 32'hfeb44683 ;
			32'h001006e4 : data_o = 32'hfea44783 ;
			32'h001006e8 : data_o = 32'h97b6078e ;
			32'h001006ec : data_o = 32'h078d078a ;
			32'h001006f0 : data_o = 32'h97221741 ;
			32'h001006f4 : data_o = 32'hec474703 ;
			32'h001006f8 : data_o = 32'h97a217c1 ;
			32'h001006fc : data_o = 32'he2e78e23 ;
			32'h00100700 : data_o = 32'hfea44783 ;
			32'h00100704 : data_o = 32'h05230785 ;
			32'h00100708 : data_o = 32'h4703fef4 ;
			32'h0010070c : data_o = 32'h478dfea4 ;
			32'h00100710 : data_o = 32'hece7fee3 ;
			32'h00100714 : data_o = 32'hfeb44783 ;
			32'h00100718 : data_o = 32'h05a30785 ;
			32'h0010071c : data_o = 32'h4703fef4 ;
			32'h00100720 : data_o = 32'h479dfeb4 ;
			32'h00100724 : data_o = 32'hece7f1e3 ;
			32'h00100728 : data_o = 32'h00001517 ;
			32'h0010072c : data_o = 32'h46c50513 ;
			32'h00100730 : data_o = 32'h151732c1 ;
			32'h00100734 : data_o = 32'h05130000 ;
			32'h00100738 : data_o = 32'h3a5d47e5 ;
			32'h0010073c : data_o = 32'h800007b7 ;
			32'h00100740 : data_o = 32'h439c0791 ;
			32'h00100744 : data_o = 32'hc3858b91 ;
			32'h00100748 : data_o = 32'h00001517 ;
			32'h0010074c : data_o = 32'h47850513 ;
			32'h00100750 : data_o = 32'h00ef3245 ;
			32'h00100754 : data_o = 32'h00ef0d70 ;
			32'h00100758 : data_o = 32'h00ef0d30 ;
			32'h0010075c : data_o = 32'h00ef0cf0 ;
			32'h00100760 : data_o = 32'h00ef0cb0 ;
			32'h00100764 : data_o = 32'h07b70c70 ;
			32'h00100768 : data_o = 32'h07918000 ;
			32'h0010076c : data_o = 32'h8b85439c ;
			32'h00100770 : data_o = 32'h1e078e63 ;
			32'h00100774 : data_o = 32'h00001517 ;
			32'h00100778 : data_o = 32'h46050513 ;
			32'h0010077c : data_o = 32'h15173a95 ;
			32'h00100780 : data_o = 32'h05130000 ;
			32'h00100784 : data_o = 32'h32ad46e5 ;
			32'h00100788 : data_o = 32'h85136789 ;
			32'h0010078c : data_o = 32'h340d7107 ;
			32'h00100790 : data_o = 32'h10ef4505 ;
			32'h00100794 : data_o = 32'h45011ae0 ;
			32'h00100798 : data_o = 32'h1c8010ef ;
			32'h0010079c : data_o = 32'hfe0401a3 ;
			32'h001007a0 : data_o = 32'h0123a835 ;
			32'h001007a4 : data_o = 32'ha00dfe04 ;
			32'h001007a8 : data_o = 32'hfe344683 ;
			32'h001007ac : data_o = 32'hfe244703 ;
			32'h001007b0 : data_o = 32'heb040793 ;
			32'h001007b4 : data_o = 32'h85ba8636 ;
			32'h001007b8 : data_o = 32'h10ef853e ;
			32'h001007bc : data_o = 32'h47831c60 ;
			32'h001007c0 : data_o = 32'h0785fe24 ;
			32'h001007c4 : data_o = 32'hfef40123 ;
			32'h001007c8 : data_o = 32'hfe244703 ;
			32'h001007cc : data_o = 32'hfde3478d ;
			32'h001007d0 : data_o = 32'h4783fce7 ;
			32'h001007d4 : data_o = 32'h0785fe34 ;
			32'h001007d8 : data_o = 32'hfef401a3 ;
			32'h001007dc : data_o = 32'hfe344703 ;
			32'h001007e0 : data_o = 32'hf0e3479d ;
			32'h001007e4 : data_o = 32'h01a3fce7 ;
			32'h001007e8 : data_o = 32'ha835fe04 ;
			32'h001007ec : data_o = 32'hfe040123 ;
			32'h001007f0 : data_o = 32'h4683a00d ;
			32'h001007f4 : data_o = 32'h4703fe34 ;
			32'h001007f8 : data_o = 32'h0793fe24 ;
			32'h001007fc : data_o = 32'h8636eac4 ;
			32'h00100800 : data_o = 32'h853e85ba ;
			32'h00100804 : data_o = 32'h17c010ef ;
			32'h00100808 : data_o = 32'hfe244783 ;
			32'h0010080c : data_o = 32'h01230785 ;
			32'h00100810 : data_o = 32'h4703fef4 ;
			32'h00100814 : data_o = 32'h478dfe24 ;
			32'h00100818 : data_o = 32'hfce7fde3 ;
			32'h0010081c : data_o = 32'hfe344783 ;
			32'h00100820 : data_o = 32'h01a30785 ;
			32'h00100824 : data_o = 32'h4703fef4 ;
			32'h00100828 : data_o = 32'h479dfe34 ;
			32'h0010082c : data_o = 32'hfce7f0e3 ;
			32'h00100830 : data_o = 32'h00001517 ;
			32'h00100834 : data_o = 32'h3c450513 ;
			32'h00100838 : data_o = 32'h67893865 ;
			32'h0010083c : data_o = 32'h71078513 ;
			32'h00100840 : data_o = 32'h45053a85 ;
			32'h00100844 : data_o = 32'h0fc010ef ;
			32'h00100848 : data_o = 32'h10ef4505 ;
			32'h0010084c : data_o = 32'h01a31160 ;
			32'h00100850 : data_o = 32'ha085fe04 ;
			32'h00100854 : data_o = 32'hfe040123 ;
			32'h00100858 : data_o = 32'h4783a099 ;
			32'h0010085c : data_o = 32'h8385fe34 ;
			32'h00100860 : data_o = 32'h0ff7f793 ;
			32'h00100864 : data_o = 32'h00279713 ;
			32'h00100868 : data_o = 32'hfe244783 ;
			32'h0010086c : data_o = 32'h971397ba ;
			32'h00100870 : data_o = 32'h47830017 ;
			32'h00100874 : data_o = 32'h8b85fe34 ;
			32'h00100878 : data_o = 32'h078a97ba ;
			32'h0010087c : data_o = 32'heb440713 ;
			32'h00100880 : data_o = 32'h468397ba ;
			32'h00100884 : data_o = 32'h4703fe34 ;
			32'h00100888 : data_o = 32'h8636fe24 ;
			32'h0010088c : data_o = 32'h853e85ba ;
			32'h00100890 : data_o = 32'h0f0010ef ;
			32'h00100894 : data_o = 32'hfe244783 ;
			32'h00100898 : data_o = 32'h01230785 ;
			32'h0010089c : data_o = 32'h4703fef4 ;
			32'h001008a0 : data_o = 32'h478dfe24 ;
			32'h001008a4 : data_o = 32'hfae7fbe3 ;
			32'h001008a8 : data_o = 32'hfe344783 ;
			32'h001008ac : data_o = 32'h01a30785 ;
			32'h001008b0 : data_o = 32'h4703fef4 ;
			32'h001008b4 : data_o = 32'h479dfe34 ;
			32'h001008b8 : data_o = 32'hf8e7fee3 ;
			32'h001008bc : data_o = 32'h00001517 ;
			32'h001008c0 : data_o = 32'h33050513 ;
			32'h001008c4 : data_o = 32'h82dff0ef ;
			32'h001008c8 : data_o = 32'h85136789 ;
			32'h001008cc : data_o = 32'h30cd7107 ;
			32'h001008d0 : data_o = 32'h10ef4501 ;
			32'h001008d4 : data_o = 32'h01a308e0 ;
			32'h001008d8 : data_o = 32'ha085fe04 ;
			32'h001008dc : data_o = 32'hfe040123 ;
			32'h001008e0 : data_o = 32'h4783a099 ;
			32'h001008e4 : data_o = 32'h8385fe34 ;
			32'h001008e8 : data_o = 32'h0ff7f793 ;
			32'h001008ec : data_o = 32'h00279713 ;
			32'h001008f0 : data_o = 32'hfe244783 ;
			32'h001008f4 : data_o = 32'h971397ba ;
			32'h001008f8 : data_o = 32'h47830017 ;
			32'h001008fc : data_o = 32'h8b85fe34 ;
			32'h00100900 : data_o = 32'h078a97ba ;
			32'h00100904 : data_o = 32'heb440713 ;
			32'h00100908 : data_o = 32'h468397ba ;
			32'h0010090c : data_o = 32'h4703fe34 ;
			32'h00100910 : data_o = 32'h8636fe24 ;
			32'h00100914 : data_o = 32'h853e85ba ;
			32'h00100918 : data_o = 32'h068010ef ;
			32'h0010091c : data_o = 32'hfe244783 ;
			32'h00100920 : data_o = 32'h01230785 ;
			32'h00100924 : data_o = 32'h4703fef4 ;
			32'h00100928 : data_o = 32'h478dfe24 ;
			32'h0010092c : data_o = 32'hfae7fbe3 ;
			32'h00100930 : data_o = 32'hfe344783 ;
			32'h00100934 : data_o = 32'h01a30785 ;
			32'h00100938 : data_o = 32'h4703fef4 ;
			32'h0010093c : data_o = 32'h479dfe34 ;
			32'h00100940 : data_o = 32'hf8e7fee3 ;
			32'h00100944 : data_o = 32'h00ef4501 ;
			32'h00100948 : data_o = 32'h15177fb0 ;
			32'h0010094c : data_o = 32'h05130000 ;
			32'h00100950 : data_o = 32'hf0ef2b25 ;
			32'h00100954 : data_o = 32'h1517f9ef ;
			32'h00100958 : data_o = 32'h05130000 ;
			32'h0010095c : data_o = 32'hf0ef2ba5 ;
			32'h00100960 : data_o = 32'h6785f92f ;
			32'h00100964 : data_o = 32'h38878513 ;
			32'h00100968 : data_o = 32'h849ff0ef ;
			32'h0010096c : data_o = 32'h00ef4501 ;
			32'h00100970 : data_o = 32'h15177d30 ;
			32'h00100974 : data_o = 32'h05130000 ;
			32'h00100978 : data_o = 32'hf0ef29e5 ;
			32'h0010097c : data_o = 32'h6785f76f ;
			32'h00100980 : data_o = 32'h38878513 ;
			32'h00100984 : data_o = 32'h82dff0ef ;
			32'h00100988 : data_o = 32'h23254501 ;
			32'h0010098c : data_o = 32'h23154505 ;
			32'h00100990 : data_o = 32'h23054509 ;
			32'h00100994 : data_o = 32'h2b31450d ;
			32'h00100998 : data_o = 32'h800007b7 ;
			32'h0010099c : data_o = 32'hc3984709 ;
			32'h001009a0 : data_o = 32'hfc042c23 ;
			32'h001009a4 : data_o = 32'hfe042223 ;
			32'h001009a8 : data_o = 32'h2783a89d ;
			32'h001009ac : data_o = 32'h853efe44 ;
			32'h001009b0 : data_o = 32'h2a23217d ;
			32'h001009b4 : data_o = 32'h2783faa4 ;
			32'h001009b8 : data_o = 32'h078afe44 ;
			32'h001009bc : data_o = 32'h97a217c1 ;
			32'h001009c0 : data_o = 32'he3c7c783 ;
			32'h001009c4 : data_o = 32'h2783873e ;
			32'h001009c8 : data_o = 32'h078afe44 ;
			32'h001009cc : data_o = 32'h17c10785 ;
			32'h001009d0 : data_o = 32'hc78397a2 ;
			32'h001009d4 : data_o = 32'h07a2e3c7 ;
			32'h001009d8 : data_o = 32'h27838f5d ;
			32'h001009dc : data_o = 32'h078afe44 ;
			32'h001009e0 : data_o = 32'h17c10789 ;
			32'h001009e4 : data_o = 32'hc78397a2 ;
			32'h001009e8 : data_o = 32'h07c2e3c7 ;
			32'h001009ec : data_o = 32'h27838f5d ;
			32'h001009f0 : data_o = 32'h078afe44 ;
			32'h001009f4 : data_o = 32'h17c1078d ;
			32'h001009f8 : data_o = 32'hc78397a2 ;
			32'h001009fc : data_o = 32'h07e2e3c7 ;
			32'h00100a00 : data_o = 32'h27838f5d ;
			32'h00100a04 : data_o = 32'h0763fb44 ;
			32'h00100a08 : data_o = 32'h278300f7 ;
			32'h00100a0c : data_o = 32'h0785fd84 ;
			32'h00100a10 : data_o = 32'hfcf42c23 ;
			32'h00100a14 : data_o = 32'hfe442783 ;
			32'h00100a18 : data_o = 32'h22230785 ;
			32'h00100a1c : data_o = 32'h2703fef4 ;
			32'h00100a20 : data_o = 32'h47fdfe44 ;
			32'h00100a24 : data_o = 32'hf8e7d3e3 ;
			32'h00100a28 : data_o = 32'h00001517 ;
			32'h00100a2c : data_o = 32'h1f050513 ;
			32'h00100a30 : data_o = 32'hec0ff0ef ;
			32'h00100a34 : data_o = 32'hfd842503 ;
			32'h00100a38 : data_o = 32'h45293c21 ;
			32'h00100a3c : data_o = 32'h6d4000ef ;
			32'h00100a40 : data_o = 32'he2042423 ;
			32'h00100a44 : data_o = 32'h00ef4505 ;
			32'h00100a48 : data_o = 32'h00ef1570 ;
			32'h00100a4c : data_o = 32'h00ef5fb0 ;
			32'h00100a50 : data_o = 32'h15176bf0 ;
			32'h00100a54 : data_o = 32'h05130000 ;
			32'h00100a58 : data_o = 32'hf0ef1be5 ;
			32'h00100a5c : data_o = 32'h6785e96f ;
			32'h00100a60 : data_o = 32'h38878513 ;
			32'h00100a64 : data_o = 32'hf4cff0ef ;
			32'h00100a68 : data_o = 32'h4b000793 ;
			32'h00100a6c : data_o = 32'hfcf42e23 ;
			32'h00100a70 : data_o = 32'h1517aa71 ;
			32'h00100a74 : data_o = 32'h05130000 ;
			32'h00100a78 : data_o = 32'hf0ef1b65 ;
			32'h00100a7c : data_o = 32'h2503e76f ;
			32'h00100a80 : data_o = 32'h3c89fdc4 ;
			32'h00100a84 : data_o = 32'h03a00513 ;
			32'h00100a88 : data_o = 32'h45292561 ;
			32'h00100a8c : data_o = 32'h05132551 ;
			32'h00100a90 : data_o = 32'hf0ef3e80 ;
			32'h00100a94 : data_o = 32'h2a23f1ef ;
			32'h00100a98 : data_o = 32'h2823fc04 ;
			32'h00100a9c : data_o = 32'h2423fc04 ;
			32'h00100aa0 : data_o = 32'h07a3fc04 ;
			32'h00100aa4 : data_o = 32'ha0edfc04 ;
			32'h00100aa8 : data_o = 32'hfc040723 ;
			32'h00100aac : data_o = 32'h06a3a8c1 ;
			32'h00100ab0 : data_o = 32'ha85dfc04 ;
			32'h00100ab4 : data_o = 32'hfc040623 ;
			32'h00100ab8 : data_o = 32'h4783a871 ;
			32'h00100abc : data_o = 32'h0423fcf4 ;
			32'h00100ac0 : data_o = 32'h4783e2f4 ;
			32'h00100ac4 : data_o = 32'h04a3fce4 ;
			32'h00100ac8 : data_o = 32'h4783e2f4 ;
			32'h00100acc : data_o = 32'h0523fcd4 ;
			32'h00100ad0 : data_o = 32'h4783e2f4 ;
			32'h00100ad4 : data_o = 32'h05a3fcc4 ;
			32'h00100ad8 : data_o = 32'h0793e2f4 ;
			32'h00100adc : data_o = 32'h853ee284 ;
			32'h00100ae0 : data_o = 32'h4cf000ef ;
			32'h00100ae4 : data_o = 32'h521000ef ;
			32'h00100ae8 : data_o = 32'h0000100f ;
			32'h00100aec : data_o = 32'h10500073 ;
			32'h00100af0 : data_o = 32'h000ff797 ;
			32'h00100af4 : data_o = 32'h51878793 ;
			32'h00100af8 : data_o = 32'h0693439c ;
			32'h00100afc : data_o = 32'h0713e284 ;
			32'h00100b00 : data_o = 32'h8636e2c4 ;
			32'h00100b04 : data_o = 32'h853e85ba ;
			32'h00100b08 : data_o = 32'hef8ff0ef ;
			32'h00100b0c : data_o = 32'h2783872a ;
			32'h00100b10 : data_o = 32'h97bafd44 ;
			32'h00100b14 : data_o = 32'hfcf42a23 ;
			32'h00100b18 : data_o = 32'h000ff797 ;
			32'h00100b1c : data_o = 32'h4f078793 ;
			32'h00100b20 : data_o = 32'h0693439c ;
			32'h00100b24 : data_o = 32'h0713e284 ;
			32'h00100b28 : data_o = 32'h8636e2c4 ;
			32'h00100b2c : data_o = 32'h853e85ba ;
			32'h00100b30 : data_o = 32'hfdcff0ef ;
			32'h00100b34 : data_o = 32'h2783872a ;
			32'h00100b38 : data_o = 32'h97bafd04 ;
			32'h00100b3c : data_o = 32'hfcf42823 ;
			32'h00100b40 : data_o = 32'hfc842783 ;
			32'h00100b44 : data_o = 32'h24230791 ;
			32'h00100b48 : data_o = 32'h4783fcf4 ;
			32'h00100b4c : data_o = 32'h0785fcc4 ;
			32'h00100b50 : data_o = 32'hfcf40623 ;
			32'h00100b54 : data_o = 32'hfcc44703 ;
			32'h00100b58 : data_o = 32'hf0e3479d ;
			32'h00100b5c : data_o = 32'h4783f6e7 ;
			32'h00100b60 : data_o = 32'h0785fcd4 ;
			32'h00100b64 : data_o = 32'hfcf406a3 ;
			32'h00100b68 : data_o = 32'hfcd44703 ;
			32'h00100b6c : data_o = 32'hf3e3479d ;
			32'h00100b70 : data_o = 32'h4783f4e7 ;
			32'h00100b74 : data_o = 32'h0785fce4 ;
			32'h00100b78 : data_o = 32'hfcf40723 ;
			32'h00100b7c : data_o = 32'hfce44703 ;
			32'h00100b80 : data_o = 32'hf6e3479d ;
			32'h00100b84 : data_o = 32'h4783f2e7 ;
			32'h00100b88 : data_o = 32'h0785fcf4 ;
			32'h00100b8c : data_o = 32'hfcf407a3 ;
			32'h00100b90 : data_o = 32'hfcf44703 ;
			32'h00100b94 : data_o = 32'hf9e3479d ;
			32'h00100b98 : data_o = 32'h4529f0e7 ;
			32'h00100b9c : data_o = 32'h15172b95 ;
			32'h00100ba0 : data_o = 32'h05130000 ;
			32'h00100ba4 : data_o = 32'hf0ef0965 ;
			32'h00100ba8 : data_o = 32'h2503d4af ;
			32'h00100bac : data_o = 32'hf0effd44 ;
			32'h00100bb0 : data_o = 32'h05138a3f ;
			32'h00100bb4 : data_o = 32'h2ba903a0 ;
			32'h00100bb8 : data_o = 32'h2b994529 ;
			32'h00100bbc : data_o = 32'h00001517 ;
			32'h00100bc0 : data_o = 32'h08450513 ;
			32'h00100bc4 : data_o = 32'hd2cff0ef ;
			32'h00100bc8 : data_o = 32'hfd042703 ;
			32'h00100bcc : data_o = 32'h0ff00793 ;
			32'h00100bd0 : data_o = 32'h02f757b3 ;
			32'h00100bd4 : data_o = 32'hf0ef853e ;
			32'h00100bd8 : data_o = 32'h051387bf ;
			32'h00100bdc : data_o = 32'h2b0d03a0 ;
			32'h00100be0 : data_o = 32'h233d4529 ;
			32'h00100be4 : data_o = 32'h00001517 ;
			32'h00100be8 : data_o = 32'h06450513 ;
			32'h00100bec : data_o = 32'hd04ff0ef ;
			32'h00100bf0 : data_o = 32'hfc842503 ;
			32'h00100bf4 : data_o = 32'h85dff0ef ;
			32'h00100bf8 : data_o = 32'h03a00513 ;
			32'h00100bfc : data_o = 32'h45292b11 ;
			32'h00100c00 : data_o = 32'h27832b01 ;
			32'h00100c04 : data_o = 32'h17d9fdc4 ;
			32'h00100c08 : data_o = 32'hfcf42e23 ;
			32'h00100c0c : data_o = 32'hfdc42703 ;
			32'h00100c10 : data_o = 32'h32000793 ;
			32'h00100c14 : data_o = 32'he4e7efe3 ;
			32'h00100c18 : data_o = 32'h32000793 ;
			32'h00100c1c : data_o = 32'hfcf42e23 ;
			32'h00100c20 : data_o = 32'h1517aa79 ;
			32'h00100c24 : data_o = 32'h05130000 ;
			32'h00100c28 : data_o = 32'hf0ef0065 ;
			32'h00100c2c : data_o = 32'h2503cc6f ;
			32'h00100c30 : data_o = 32'hf0effdc4 ;
			32'h00100c34 : data_o = 32'h05138a3f ;
			32'h00100c38 : data_o = 32'h29d903a0 ;
			32'h00100c3c : data_o = 32'h29c94529 ;
			32'h00100c40 : data_o = 32'h3e800513 ;
			32'h00100c44 : data_o = 32'hd6cff0ef ;
			32'h00100c48 : data_o = 32'hfc042223 ;
			32'h00100c4c : data_o = 32'hfc042023 ;
			32'h00100c50 : data_o = 32'hfa042c23 ;
			32'h00100c54 : data_o = 32'hfa040fa3 ;
			32'h00100c58 : data_o = 32'h0f23a0ed ;
			32'h00100c5c : data_o = 32'ha8c1fa04 ;
			32'h00100c60 : data_o = 32'hfa040ea3 ;
			32'h00100c64 : data_o = 32'h0e23a85d ;
			32'h00100c68 : data_o = 32'ha871fa04 ;
			32'h00100c6c : data_o = 32'hfbf44783 ;
			32'h00100c70 : data_o = 32'he2f40423 ;
			32'h00100c74 : data_o = 32'hfbe44783 ;
			32'h00100c78 : data_o = 32'he2f404a3 ;
			32'h00100c7c : data_o = 32'hfbd44783 ;
			32'h00100c80 : data_o = 32'he2f40523 ;
			32'h00100c84 : data_o = 32'hfbc44783 ;
			32'h00100c88 : data_o = 32'he2f405a3 ;
			32'h00100c8c : data_o = 32'he2840793 ;
			32'h00100c90 : data_o = 32'h00ef853e ;
			32'h00100c94 : data_o = 32'h00ef31d0 ;
			32'h00100c98 : data_o = 32'h100f36f0 ;
			32'h00100c9c : data_o = 32'h00730000 ;
			32'h00100ca0 : data_o = 32'hf7971050 ;
			32'h00100ca4 : data_o = 32'h8793000f ;
			32'h00100ca8 : data_o = 32'h439c3667 ;
			32'h00100cac : data_o = 32'he2840693 ;
			32'h00100cb0 : data_o = 32'he2c40713 ;
			32'h00100cb4 : data_o = 32'h85ba8636 ;
			32'h00100cb8 : data_o = 32'hf0ef853e ;
			32'h00100cbc : data_o = 32'h872ad46f ;
			32'h00100cc0 : data_o = 32'hfc442783 ;
			32'h00100cc4 : data_o = 32'h222397ba ;
			32'h00100cc8 : data_o = 32'hf797fcf4 ;
			32'h00100ccc : data_o = 32'h8793000f ;
			32'h00100cd0 : data_o = 32'h439c33e7 ;
			32'h00100cd4 : data_o = 32'he2840693 ;
			32'h00100cd8 : data_o = 32'he2c40713 ;
			32'h00100cdc : data_o = 32'h85ba8636 ;
			32'h00100ce0 : data_o = 32'hf0ef853e ;
			32'h00100ce4 : data_o = 32'h872ae2af ;
			32'h00100ce8 : data_o = 32'hfc042783 ;
			32'h00100cec : data_o = 32'h202397ba ;
			32'h00100cf0 : data_o = 32'h2783fcf4 ;
			32'h00100cf4 : data_o = 32'h0791fb84 ;
			32'h00100cf8 : data_o = 32'hfaf42c23 ;
			32'h00100cfc : data_o = 32'hfbc44783 ;
			32'h00100d00 : data_o = 32'h0e230785 ;
			32'h00100d04 : data_o = 32'h4703faf4 ;
			32'h00100d08 : data_o = 32'h479dfbc4 ;
			32'h00100d0c : data_o = 32'hf6e7f0e3 ;
			32'h00100d10 : data_o = 32'hfbd44783 ;
			32'h00100d14 : data_o = 32'h0ea30785 ;
			32'h00100d18 : data_o = 32'h4703faf4 ;
			32'h00100d1c : data_o = 32'h479dfbd4 ;
			32'h00100d20 : data_o = 32'hf4e7f3e3 ;
			32'h00100d24 : data_o = 32'hfbe44783 ;
			32'h00100d28 : data_o = 32'h0f230785 ;
			32'h00100d2c : data_o = 32'h4703faf4 ;
			32'h00100d30 : data_o = 32'h479dfbe4 ;
			32'h00100d34 : data_o = 32'hf2e7f6e3 ;
			32'h00100d38 : data_o = 32'hfbf44783 ;
			32'h00100d3c : data_o = 32'h0fa30785 ;
			32'h00100d40 : data_o = 32'h4703faf4 ;
			32'h00100d44 : data_o = 32'h479dfbf4 ;
			32'h00100d48 : data_o = 32'hf0e7f9e3 ;
			32'h00100d4c : data_o = 32'h26c94529 ;
			32'h00100d50 : data_o = 32'h00001517 ;
			32'h00100d54 : data_o = 32'hee450513 ;
			32'h00100d58 : data_o = 32'hb98ff0ef ;
			32'h00100d5c : data_o = 32'hfc442503 ;
			32'h00100d60 : data_o = 32'hef0ff0ef ;
			32'h00100d64 : data_o = 32'h03a00513 ;
			32'h00100d68 : data_o = 32'h45292665 ;
			32'h00100d6c : data_o = 32'h15172655 ;
			32'h00100d70 : data_o = 32'h05130000 ;
			32'h00100d74 : data_o = 32'hf0efed25 ;
			32'h00100d78 : data_o = 32'h2703b7af ;
			32'h00100d7c : data_o = 32'h0793fc04 ;
			32'h00100d80 : data_o = 32'h57b30ff0 ;
			32'h00100d84 : data_o = 32'h853e02f7 ;
			32'h00100d88 : data_o = 32'hec8ff0ef ;
			32'h00100d8c : data_o = 32'h03a00513 ;
			32'h00100d90 : data_o = 32'h45292641 ;
			32'h00100d94 : data_o = 32'h15172eb5 ;
			32'h00100d98 : data_o = 32'h05130000 ;
			32'h00100d9c : data_o = 32'hf0efeb25 ;
			32'h00100da0 : data_o = 32'h2503b52f ;
			32'h00100da4 : data_o = 32'hf0effb84 ;
			32'h00100da8 : data_o = 32'h0513eaaf ;
			32'h00100dac : data_o = 32'h268d03a0 ;
			32'h00100db0 : data_o = 32'h2eb94529 ;
			32'h00100db4 : data_o = 32'hfdc42783 ;
			32'h00100db8 : data_o = 32'h2e2317ed ;
			32'h00100dbc : data_o = 32'h2703fcf4 ;
			32'h00100dc0 : data_o = 32'h0793fdc4 ;
			32'h00100dc4 : data_o = 32'heee32580 ;
			32'h00100dc8 : data_o = 32'h1517e4e7 ;
			32'h00100dcc : data_o = 32'h05130000 ;
			32'h00100dd0 : data_o = 32'hf0efe8a5 ;
			32'h00100dd4 : data_o = 32'h4781b1ef ;
			32'h00100dd8 : data_o = 32'h2083853e ;
			32'h00100ddc : data_o = 32'h24031dc1 ;
			32'h00100de0 : data_o = 32'h613d1d81 ;
			32'h00100de4 : data_o = 32'h71798082 ;
			32'h00100de8 : data_o = 32'h1800d622 ;
			32'h00100dec : data_o = 32'hfca42e23 ;
			32'h00100df0 : data_o = 32'hfcb42c23 ;
			32'h00100df4 : data_o = 32'hfe042623 ;
			32'h00100df8 : data_o = 32'h477da0a1 ;
			32'h00100dfc : data_o = 32'hfec42783 ;
			32'h00100e00 : data_o = 32'h40f707b3 ;
			32'h00100e04 : data_o = 32'hfdc42703 ;
			32'h00100e08 : data_o = 32'h00f757b3 ;
			32'h00100e0c : data_o = 32'hcb998b85 ;
			32'h00100e10 : data_o = 32'hfec42783 ;
			32'h00100e14 : data_o = 32'hfd842703 ;
			32'h00100e18 : data_o = 32'h071397ba ;
			32'h00100e1c : data_o = 32'h80230310 ;
			32'h00100e20 : data_o = 32'ha81100e7 ;
			32'h00100e24 : data_o = 32'hfec42783 ;
			32'h00100e28 : data_o = 32'hfd842703 ;
			32'h00100e2c : data_o = 32'h071397ba ;
			32'h00100e30 : data_o = 32'h80230300 ;
			32'h00100e34 : data_o = 32'h278300e7 ;
			32'h00100e38 : data_o = 32'h0785fec4 ;
			32'h00100e3c : data_o = 32'hfef42623 ;
			32'h00100e40 : data_o = 32'hfec42703 ;
			32'h00100e44 : data_o = 32'hdae347fd ;
			32'h00100e48 : data_o = 32'h2783fae7 ;
			32'h00100e4c : data_o = 32'h8793fd84 ;
			32'h00100e50 : data_o = 32'h80230207 ;
			32'h00100e54 : data_o = 32'h00010007 ;
			32'h00100e58 : data_o = 32'h61455432 ;
			32'h00100e5c : data_o = 32'h11018082 ;
			32'h00100e60 : data_o = 32'h1000ce22 ;
			32'h00100e64 : data_o = 32'hfea42623 ;
			32'h00100e68 : data_o = 32'hfec42703 ;
			32'h00100e6c : data_o = 32'h1c0007b7 ;
			32'h00100e70 : data_o = 32'h20078793 ;
			32'h00100e74 : data_o = 32'h078a97ba ;
			32'h00100e78 : data_o = 32'h853e439c ;
			32'h00100e7c : data_o = 32'h61054472 ;
			32'h00100e80 : data_o = 32'h11018082 ;
			32'h00100e84 : data_o = 32'h1000ce22 ;
			32'h00100e88 : data_o = 32'hfea42623 ;
			32'h00100e8c : data_o = 32'hfeb42423 ;
			32'h00100e90 : data_o = 32'hfe842783 ;
			32'h00100e94 : data_o = 32'hfec42703 ;
			32'h00100e98 : data_o = 32'h00f757b3 ;
			32'h00100e9c : data_o = 32'hc7818b85 ;
			32'h00100ea0 : data_o = 32'h03100793 ;
			32'h00100ea4 : data_o = 32'h0793a019 ;
			32'h00100ea8 : data_o = 32'h853e0300 ;
			32'h00100eac : data_o = 32'h61054472 ;
			32'h00100eb0 : data_o = 32'h715d8082 ;
			32'h00100eb4 : data_o = 32'hc4a2c686 ;
			32'h00100eb8 : data_o = 32'h0880c2a6 ;
			32'h00100ebc : data_o = 32'hfaa42e23 ;
			32'h00100ec0 : data_o = 32'hfbc42703 ;
			32'h00100ec4 : data_o = 32'hf463478d ;
			32'h00100ec8 : data_o = 32'h000100e7 ;
			32'h00100ecc : data_o = 32'h2623aa81 ;
			32'h00100ed0 : data_o = 32'ha0a5fe04 ;
			32'h00100ed4 : data_o = 32'hfec42783 ;
			32'h00100ed8 : data_o = 32'h00279713 ;
			32'h00100edc : data_o = 32'hfbc42783 ;
			32'h00100ee0 : data_o = 32'h971397ba ;
			32'h00100ee4 : data_o = 32'h27830017 ;
			32'h00100ee8 : data_o = 32'h9493fec4 ;
			32'h00100eec : data_o = 32'h853a0017 ;
			32'h00100ef0 : data_o = 32'h872a37bd ;
			32'h00100ef4 : data_o = 32'h00249793 ;
			32'h00100ef8 : data_o = 32'h97a217c1 ;
			32'h00100efc : data_o = 32'hfce7a823 ;
			32'h00100f00 : data_o = 32'hfec42783 ;
			32'h00100f04 : data_o = 32'h00279713 ;
			32'h00100f08 : data_o = 32'hfbc42783 ;
			32'h00100f0c : data_o = 32'h078697ba ;
			32'h00100f10 : data_o = 32'h00178713 ;
			32'h00100f14 : data_o = 32'hfec42783 ;
			32'h00100f18 : data_o = 32'h84930786 ;
			32'h00100f1c : data_o = 32'h853a0017 ;
			32'h00100f20 : data_o = 32'h872a3f3d ;
			32'h00100f24 : data_o = 32'h00249793 ;
			32'h00100f28 : data_o = 32'h97a217c1 ;
			32'h00100f2c : data_o = 32'hfce7a823 ;
			32'h00100f30 : data_o = 32'hfec42783 ;
			32'h00100f34 : data_o = 32'h26230785 ;
			32'h00100f38 : data_o = 32'h2703fef4 ;
			32'h00100f3c : data_o = 32'h478dfec4 ;
			32'h00100f40 : data_o = 32'hf8e7fae3 ;
			32'h00100f44 : data_o = 32'h22e94529 ;
			32'h00100f48 : data_o = 32'hfe042223 ;
			32'h00100f4c : data_o = 32'h2423a0c9 ;
			32'h00100f50 : data_o = 32'ha055fe04 ;
			32'h00100f54 : data_o = 32'h07c00513 ;
			32'h00100f58 : data_o = 32'h20232a65 ;
			32'h00100f5c : data_o = 32'ha8bdfe04 ;
			32'h00100f60 : data_o = 32'hfe442703 ;
			32'h00100f64 : data_o = 32'hca63478d ;
			32'h00100f68 : data_o = 32'h278302e7 ;
			32'h00100f6c : data_o = 32'h0786fe84 ;
			32'h00100f70 : data_o = 32'h17c1078a ;
			32'h00100f74 : data_o = 32'ha68397a2 ;
			32'h00100f78 : data_o = 32'h2783fd07 ;
			32'h00100f7c : data_o = 32'h078efe44 ;
			32'h00100f80 : data_o = 32'h00778713 ;
			32'h00100f84 : data_o = 32'hfe042783 ;
			32'h00100f88 : data_o = 32'h40f707b3 ;
			32'h00100f8c : data_o = 32'h853685be ;
			32'h00100f90 : data_o = 32'h87aa3dcd ;
			32'h00100f94 : data_o = 32'h2aad853e ;
			32'h00100f98 : data_o = 32'h2783a815 ;
			32'h00100f9c : data_o = 32'h0786fe84 ;
			32'h00100fa0 : data_o = 32'h078a0785 ;
			32'h00100fa4 : data_o = 32'h97a217c1 ;
			32'h00100fa8 : data_o = 32'hfd07a683 ;
			32'h00100fac : data_o = 32'hfe442783 ;
			32'h00100fb0 : data_o = 32'h078e17f1 ;
			32'h00100fb4 : data_o = 32'h00778713 ;
			32'h00100fb8 : data_o = 32'hfe042783 ;
			32'h00100fbc : data_o = 32'h40f707b3 ;
			32'h00100fc0 : data_o = 32'h853685be ;
			32'h00100fc4 : data_o = 32'h87aa3d7d ;
			32'h00100fc8 : data_o = 32'h2299853e ;
			32'h00100fcc : data_o = 32'h07c00513 ;
			32'h00100fd0 : data_o = 32'h27832281 ;
			32'h00100fd4 : data_o = 32'h0785fe04 ;
			32'h00100fd8 : data_o = 32'hfef42023 ;
			32'h00100fdc : data_o = 32'hfe042703 ;
			32'h00100fe0 : data_o = 32'hdfe3479d ;
			32'h00100fe4 : data_o = 32'h0513f6e7 ;
			32'h00100fe8 : data_o = 32'h221d0200 ;
			32'h00100fec : data_o = 32'hfe842783 ;
			32'h00100ff0 : data_o = 32'h24230785 ;
			32'h00100ff4 : data_o = 32'h2703fef4 ;
			32'h00100ff8 : data_o = 32'h478dfe84 ;
			32'h00100ffc : data_o = 32'hf4e7dce3 ;
			32'h00101000 : data_o = 32'h22394529 ;
			32'h00101004 : data_o = 32'hfe442783 ;
			32'h00101008 : data_o = 32'h22230785 ;
			32'h0010100c : data_o = 32'h2703fef4 ;
			32'h00101010 : data_o = 32'h479dfe44 ;
			32'h00101014 : data_o = 32'hf2e7dde3 ;
			32'h00101018 : data_o = 32'h28dd4529 ;
			32'h0010101c : data_o = 32'h40b60001 ;
			32'h00101020 : data_o = 32'h44964426 ;
			32'h00101024 : data_o = 32'h80826161 ;
			32'h00101028 : data_o = 32'hce061101 ;
			32'h0010102c : data_o = 32'h1000cc22 ;
			32'h00101030 : data_o = 32'hfe042223 ;
			32'h00101034 : data_o = 32'h202357fd ;
			32'h00101038 : data_o = 32'h1517fef4 ;
			32'h0010103c : data_o = 32'h05130000 ;
			32'h00101040 : data_o = 32'hf0efca25 ;
			32'h00101044 : data_o = 32'h67858aef ;
			32'h00101048 : data_o = 32'h38878513 ;
			32'h0010104c : data_o = 32'h964ff0ef ;
			32'h00101050 : data_o = 32'h00ef4505 ;
			32'h00101054 : data_o = 32'h45050ef0 ;
			32'h00101058 : data_o = 32'h109000ef ;
			32'h0010105c : data_o = 32'hfe042623 ;
			32'h00101060 : data_o = 32'h2423a091 ;
			32'h00101064 : data_o = 32'ha02dfe04 ;
			32'h00101068 : data_o = 32'hfe842783 ;
			32'h0010106c : data_o = 32'h0ff7f713 ;
			32'h00101070 : data_o = 32'hfec42783 ;
			32'h00101074 : data_o = 32'h0ff7f693 ;
			32'h00101078 : data_o = 32'hfe440793 ;
			32'h0010107c : data_o = 32'h85ba8636 ;
			32'h00101080 : data_o = 32'h00ef853e ;
			32'h00101084 : data_o = 32'h27830ff0 ;
			32'h00101088 : data_o = 32'h0785fe84 ;
			32'h0010108c : data_o = 32'hfef42423 ;
			32'h00101090 : data_o = 32'hfe842703 ;
			32'h00101094 : data_o = 32'hd9e3478d ;
			32'h00101098 : data_o = 32'h2783fce7 ;
			32'h0010109c : data_o = 32'h0785fec4 ;
			32'h001010a0 : data_o = 32'hfef42623 ;
			32'h001010a4 : data_o = 32'hfec42703 ;
			32'h001010a8 : data_o = 32'hdce3479d ;
			32'h001010ac : data_o = 32'h2623fae7 ;
			32'h001010b0 : data_o = 32'ha091fe04 ;
			32'h001010b4 : data_o = 32'hfe042423 ;
			32'h001010b8 : data_o = 32'h2783a02d ;
			32'h001010bc : data_o = 32'hf713fe84 ;
			32'h001010c0 : data_o = 32'h27830ff7 ;
			32'h001010c4 : data_o = 32'hf693fec4 ;
			32'h001010c8 : data_o = 32'h07930ff7 ;
			32'h001010cc : data_o = 32'h8636fe04 ;
			32'h001010d0 : data_o = 32'h853e85ba ;
			32'h001010d4 : data_o = 32'h0ad000ef ;
			32'h001010d8 : data_o = 32'hfe842783 ;
			32'h001010dc : data_o = 32'h24230785 ;
			32'h001010e0 : data_o = 32'h2703fef4 ;
			32'h001010e4 : data_o = 32'h478dfe84 ;
			32'h001010e8 : data_o = 32'hfce7d9e3 ;
			32'h001010ec : data_o = 32'hfec42783 ;
			32'h001010f0 : data_o = 32'h26230785 ;
			32'h001010f4 : data_o = 32'h2703fef4 ;
			32'h001010f8 : data_o = 32'h479dfec4 ;
			32'h001010fc : data_o = 32'hfae7dce3 ;
			32'h00101100 : data_o = 32'h00ef4501 ;
			32'h00101104 : data_o = 32'h000103f0 ;
			32'h00101108 : data_o = 32'h446240f2 ;
			32'h0010110c : data_o = 32'h80826105 ;
			32'h00101110 : data_o = 32'hce061101 ;
			32'h00101114 : data_o = 32'h1000cc22 ;
			32'h00101118 : data_o = 32'h07a387aa ;
			32'h0010111c : data_o = 32'h4703fef4 ;
			32'h00101120 : data_o = 32'h47a9fef4 ;
			32'h00101124 : data_o = 32'h00f71663 ;
			32'h00101128 : data_o = 32'h153745b5 ;
			32'h0010112c : data_o = 32'h2e2d8000 ;
			32'h00101130 : data_o = 32'hfef44783 ;
			32'h00101134 : data_o = 32'h153785be ;
			32'h00101138 : data_o = 32'h263d8000 ;
			32'h0010113c : data_o = 32'hfef44783 ;
			32'h00101140 : data_o = 32'h40f2853e ;
			32'h00101144 : data_o = 32'h61054462 ;
			32'h00101148 : data_o = 32'h11418082 ;
			32'h0010114c : data_o = 32'hc422c606 ;
			32'h00101150 : data_o = 32'h15370800 ;
			32'h00101154 : data_o = 32'h24c58000 ;
			32'h00101158 : data_o = 32'h853e87aa ;
			32'h0010115c : data_o = 32'h442240b2 ;
			32'h00101160 : data_o = 32'h80820141 ;
			32'h00101164 : data_o = 32'hce061101 ;
			32'h00101168 : data_o = 32'h1000cc22 ;
			32'h0010116c : data_o = 32'hfea42623 ;
			32'h00101170 : data_o = 32'h2783a819 ;
			32'h00101174 : data_o = 32'h8713fec4 ;
			32'h00101178 : data_o = 32'h26230017 ;
			32'h0010117c : data_o = 32'hc783fee4 ;
			32'h00101180 : data_o = 32'h853e0007 ;
			32'h00101184 : data_o = 32'h27833771 ;
			32'h00101188 : data_o = 32'hc783fec4 ;
			32'h0010118c : data_o = 32'hf3f50007 ;
			32'h00101190 : data_o = 32'h853e4781 ;
			32'h00101194 : data_o = 32'h446240f2 ;
			32'h00101198 : data_o = 32'h80826105 ;
			32'h0010119c : data_o = 32'hd6067179 ;
			32'h001011a0 : data_o = 32'h1800d422 ;
			32'h001011a4 : data_o = 32'hfca42e23 ;
			32'h001011a8 : data_o = 32'hfe042623 ;
			32'h001011ac : data_o = 32'h2783a891 ;
			32'h001011b0 : data_o = 32'h83f1fdc4 ;
			32'h001011b4 : data_o = 32'hfef42423 ;
			32'h001011b8 : data_o = 32'hfe842703 ;
			32'h001011bc : data_o = 32'hcd6347a5 ;
			32'h001011c0 : data_o = 32'h278300e7 ;
			32'h001011c4 : data_o = 32'hf793fe84 ;
			32'h001011c8 : data_o = 32'h87930ff7 ;
			32'h001011cc : data_o = 32'hf7930307 ;
			32'h001011d0 : data_o = 32'h853e0ff7 ;
			32'h001011d4 : data_o = 32'ha8193f35 ;
			32'h001011d8 : data_o = 32'hfe842783 ;
			32'h001011dc : data_o = 32'h0ff7f793 ;
			32'h001011e0 : data_o = 32'h03778793 ;
			32'h001011e4 : data_o = 32'h0ff7f793 ;
			32'h001011e8 : data_o = 32'h371d853e ;
			32'h001011ec : data_o = 32'hfdc42783 ;
			32'h001011f0 : data_o = 32'h2e230792 ;
			32'h001011f4 : data_o = 32'h2783fcf4 ;
			32'h001011f8 : data_o = 32'h0785fec4 ;
			32'h001011fc : data_o = 32'hfef42623 ;
			32'h00101200 : data_o = 32'hfec42703 ;
			32'h00101204 : data_o = 32'hd4e3479d ;
			32'h00101208 : data_o = 32'h0001fae7 ;
			32'h0010120c : data_o = 32'h50b20001 ;
			32'h00101210 : data_o = 32'h61455422 ;
			32'h00101214 : data_o = 32'h11418082 ;
			32'h00101218 : data_o = 32'h0800c622 ;
			32'h0010121c : data_o = 32'h000207b7 ;
			32'h00101220 : data_o = 32'h470507a1 ;
			32'h00101224 : data_o = 32'h0001c398 ;
			32'h00101228 : data_o = 32'h01414432 ;
			32'h0010122c : data_o = 32'h11018082 ;
			32'h00101230 : data_o = 32'h1000ce22 ;
			32'h00101234 : data_o = 32'h341027f3 ;
			32'h00101238 : data_o = 32'hfef42623 ;
			32'h0010123c : data_o = 32'hfec42783 ;
			32'h00101240 : data_o = 32'h4472853e ;
			32'h00101244 : data_o = 32'h80826105 ;
			32'h00101248 : data_o = 32'hce221101 ;
			32'h0010124c : data_o = 32'h27f31000 ;
			32'h00101250 : data_o = 32'h26233420 ;
			32'h00101254 : data_o = 32'h2783fef4 ;
			32'h00101258 : data_o = 32'h853efec4 ;
			32'h0010125c : data_o = 32'h61054472 ;
			32'h00101260 : data_o = 32'h11018082 ;
			32'h00101264 : data_o = 32'h1000ce22 ;
			32'h00101268 : data_o = 32'h343027f3 ;
			32'h0010126c : data_o = 32'hfef42623 ;
			32'h00101270 : data_o = 32'hfec42783 ;
			32'h00101274 : data_o = 32'h4472853e ;
			32'h00101278 : data_o = 32'h80826105 ;
			32'h0010127c : data_o = 32'hce221101 ;
			32'h00101280 : data_o = 32'h27f31000 ;
			32'h00101284 : data_o = 32'h2623b000 ;
			32'h00101288 : data_o = 32'h2783fef4 ;
			32'h0010128c : data_o = 32'h853efec4 ;
			32'h00101290 : data_o = 32'h61054472 ;
			32'h00101294 : data_o = 32'h11418082 ;
			32'h00101298 : data_o = 32'h0800c622 ;
			32'h0010129c : data_o = 32'hb0001073 ;
			32'h001012a0 : data_o = 32'h44320001 ;
			32'h001012a4 : data_o = 32'h80820141 ;
			32'h001012a8 : data_o = 32'hd6227179 ;
			32'h001012ac : data_o = 32'h2e231800 ;
			32'h001012b0 : data_o = 32'h2c23fca4 ;
			32'h001012b4 : data_o = 32'h2703fcb4 ;
			32'h001012b8 : data_o = 32'h47fdfdc4 ;
			32'h001012bc : data_o = 32'h00e7f463 ;
			32'h001012c0 : data_o = 32'ha8794785 ;
			32'h001012c4 : data_o = 32'h000ff797 ;
			32'h001012c8 : data_o = 32'hd3c78793 ;
			32'h001012cc : data_o = 32'h27834398 ;
			32'h001012d0 : data_o = 32'h078afdc4 ;
			32'h001012d4 : data_o = 32'h262397ba ;
			32'h001012d8 : data_o = 32'h2703fef4 ;
			32'h001012dc : data_o = 32'h2783fd84 ;
			32'h001012e0 : data_o = 32'h07b3fec4 ;
			32'h001012e4 : data_o = 32'h242340f7 ;
			32'h001012e8 : data_o = 32'h2703fef4 ;
			32'h001012ec : data_o = 32'h07b7fe84 ;
			32'h001012f0 : data_o = 32'h58630008 ;
			32'h001012f4 : data_o = 32'h270300f7 ;
			32'h001012f8 : data_o = 32'h07b7fe84 ;
			32'h001012fc : data_o = 32'h5463fff8 ;
			32'h00101300 : data_o = 32'h478900f7 ;
			32'h00101304 : data_o = 32'h2783a8b1 ;
			32'h00101308 : data_o = 32'h2223fe84 ;
			32'h0010130c : data_o = 32'h2783fef4 ;
			32'h00101310 : data_o = 32'h9713fe44 ;
			32'h00101314 : data_o = 32'h07b70147 ;
			32'h00101318 : data_o = 32'h8f7d7fe0 ;
			32'h0010131c : data_o = 32'hfe442783 ;
			32'h00101320 : data_o = 32'h00979693 ;
			32'h00101324 : data_o = 32'h001007b7 ;
			32'h00101328 : data_o = 32'h8f5d8ff5 ;
			32'h0010132c : data_o = 32'hfe442683 ;
			32'h00101330 : data_o = 32'h000ff7b7 ;
			32'h00101334 : data_o = 32'h8f5d8ff5 ;
			32'h00101338 : data_o = 32'hfe442783 ;
			32'h0010133c : data_o = 32'h00b79693 ;
			32'h00101340 : data_o = 32'h800007b7 ;
			32'h00101344 : data_o = 32'h8fd98ff5 ;
			32'h00101348 : data_o = 32'h06f7e793 ;
			32'h0010134c : data_o = 32'hfef42023 ;
			32'h00101350 : data_o = 32'hfec42783 ;
			32'h00101354 : data_o = 32'hfe042703 ;
			32'h00101358 : data_o = 32'h100fc398 ;
			32'h0010135c : data_o = 32'h47810000 ;
			32'h00101360 : data_o = 32'h5432853e ;
			32'h00101364 : data_o = 32'h80826145 ;
			32'h00101368 : data_o = 32'hce221101 ;
			32'h0010136c : data_o = 32'h26231000 ;
			32'h00101370 : data_o = 32'h2783fea4 ;
			32'h00101374 : data_o = 32'ha073fec4 ;
			32'h00101378 : data_o = 32'h00013047 ;
			32'h0010137c : data_o = 32'h61054472 ;
			32'h00101380 : data_o = 32'h11018082 ;
			32'h00101384 : data_o = 32'h1000ce22 ;
			32'h00101388 : data_o = 32'hfea42623 ;
			32'h0010138c : data_o = 32'hfec42783 ;
			32'h00101390 : data_o = 32'h3047b073 ;
			32'h00101394 : data_o = 32'h44720001 ;
			32'h00101398 : data_o = 32'h80826105 ;
			32'h0010139c : data_o = 32'hce221101 ;
			32'h001013a0 : data_o = 32'h26231000 ;
			32'h001013a4 : data_o = 32'h2783fea4 ;
			32'h001013a8 : data_o = 32'hc789fec4 ;
			32'h001013ac : data_o = 32'ha07347a1 ;
			32'h001013b0 : data_o = 32'ha0213007 ;
			32'h001013b4 : data_o = 32'hb07347a1 ;
			32'h001013b8 : data_o = 32'h00013007 ;
			32'h001013bc : data_o = 32'h61054472 ;
			32'h001013c0 : data_o = 32'h11418082 ;
			32'h001013c4 : data_o = 32'hc422c606 ;
			32'h001013c8 : data_o = 32'h15170800 ;
			32'h001013cc : data_o = 32'h05130000 ;
			32'h001013d0 : data_o = 32'h3b4991a5 ;
			32'h001013d4 : data_o = 32'h00001517 ;
			32'h001013d8 : data_o = 32'h92050513 ;
			32'h001013dc : data_o = 32'h15173361 ;
			32'h001013e0 : data_o = 32'h05130000 ;
			32'h001013e4 : data_o = 32'h3bbd9265 ;
			32'h001013e8 : data_o = 32'h87aa3599 ;
			32'h001013ec : data_o = 32'h337d853e ;
			32'h001013f0 : data_o = 32'h00001517 ;
			32'h001013f4 : data_o = 32'h92050513 ;
			32'h001013f8 : data_o = 32'h35b933b5 ;
			32'h001013fc : data_o = 32'h853e87aa ;
			32'h00101400 : data_o = 32'h15173b71 ;
			32'h00101404 : data_o = 32'h05130000 ;
			32'h00101408 : data_o = 32'h3ba991a5 ;
			32'h0010140c : data_o = 32'h87aa3d99 ;
			32'h00101410 : data_o = 32'h3369853e ;
			32'h00101414 : data_o = 32'h39ed4529 ;
			32'h00101418 : data_o = 32'hbffd0001 ;
			32'h0010141c : data_o = 32'hc6061141 ;
			32'h00101420 : data_o = 32'h0800c422 ;
			32'h00101424 : data_o = 32'h37896541 ;
			32'h00101428 : data_o = 32'h3f8d4505 ;
			32'h0010142c : data_o = 32'h40b20001 ;
			32'h00101430 : data_o = 32'h01414422 ;
			32'h00101434 : data_o = 32'h71798082 ;
			32'h00101438 : data_o = 32'h1800d622 ;
			32'h0010143c : data_o = 32'hfca42e23 ;
			32'h00101440 : data_o = 32'h262357fd ;
			32'h00101444 : data_o = 32'h2783fef4 ;
			32'h00101448 : data_o = 32'h07a1fdc4 ;
			32'h0010144c : data_o = 32'h8b85439c ;
			32'h00101450 : data_o = 32'h2783e791 ;
			32'h00101454 : data_o = 32'h439cfdc4 ;
			32'h00101458 : data_o = 32'hfef42623 ;
			32'h0010145c : data_o = 32'hfec42783 ;
			32'h00101460 : data_o = 32'h5432853e ;
			32'h00101464 : data_o = 32'h80826145 ;
			32'h00101468 : data_o = 32'hce221101 ;
			32'h0010146c : data_o = 32'h26231000 ;
			32'h00101470 : data_o = 32'h87aefea4 ;
			32'h00101474 : data_o = 32'hfef405a3 ;
			32'h00101478 : data_o = 32'h27830001 ;
			32'h0010147c : data_o = 32'h07a1fec4 ;
			32'h00101480 : data_o = 32'h8b89439c ;
			32'h00101484 : data_o = 32'h2783fbfd ;
			32'h00101488 : data_o = 32'h0791fec4 ;
			32'h0010148c : data_o = 32'hfeb44703 ;
			32'h00101490 : data_o = 32'h0001c398 ;
			32'h00101494 : data_o = 32'h61054472 ;
			32'h00101498 : data_o = 32'h11018082 ;
			32'h0010149c : data_o = 32'h1000ce22 ;
			32'h001014a0 : data_o = 32'hfea42423 ;
			32'h001014a4 : data_o = 32'hfeb42623 ;
			32'h001014a8 : data_o = 32'h080026b7 ;
			32'h001014ac : data_o = 32'h567d06a1 ;
			32'h001014b0 : data_o = 32'h2683c290 ;
			32'h001014b4 : data_o = 32'hd713fec4 ;
			32'h001014b8 : data_o = 32'h47810006 ;
			32'h001014bc : data_o = 32'h080026b7 ;
			32'h001014c0 : data_o = 32'h87ba06b1 ;
			32'h001014c4 : data_o = 32'h27b7c29c ;
			32'h001014c8 : data_o = 32'h07a10800 ;
			32'h001014cc : data_o = 32'hfe842703 ;
			32'h001014d0 : data_o = 32'h0001c398 ;
			32'h001014d4 : data_o = 32'h61054472 ;
			32'h001014d8 : data_o = 32'h71798082 ;
			32'h001014dc : data_o = 32'hd422d606 ;
			32'h001014e0 : data_o = 32'h2c231800 ;
			32'h001014e4 : data_o = 32'h2e23fca4 ;
			32'h001014e8 : data_o = 32'h20fdfcb4 ;
			32'h001014ec : data_o = 32'hfea42423 ;
			32'h001014f0 : data_o = 32'hfeb42623 ;
			32'h001014f4 : data_o = 32'hfe842603 ;
			32'h001014f8 : data_o = 32'hfec42683 ;
			32'h001014fc : data_o = 32'hfd842503 ;
			32'h00101500 : data_o = 32'hfdc42583 ;
			32'h00101504 : data_o = 32'h00a60733 ;
			32'h00101508 : data_o = 32'h3833883a ;
			32'h0010150c : data_o = 32'h87b300c8 ;
			32'h00101510 : data_o = 32'h06b300b6 ;
			32'h00101514 : data_o = 32'h87b600f8 ;
			32'h00101518 : data_o = 32'hfee42423 ;
			32'h0010151c : data_o = 32'hfef42623 ;
			32'h00101520 : data_o = 32'hfe842503 ;
			32'h00101524 : data_o = 32'hfec42583 ;
			32'h00101528 : data_o = 32'h00013f8d ;
			32'h0010152c : data_o = 32'h542250b2 ;
			32'h00101530 : data_o = 32'h80826145 ;
			32'h00101534 : data_o = 32'hc686715d ;
			32'h00101538 : data_o = 32'hc29ac496 ;
			32'h0010153c : data_o = 32'hde22c09e ;
			32'h00101540 : data_o = 32'hda2edc2a ;
			32'h00101544 : data_o = 32'hd636d832 ;
			32'h00101548 : data_o = 32'hd23ed43a ;
			32'h0010154c : data_o = 32'hce46d042 ;
			32'h00101550 : data_o = 32'hca76cc72 ;
			32'h00101554 : data_o = 32'hc67ec87a ;
			32'h00101558 : data_o = 32'hf7970880 ;
			32'h0010155c : data_o = 32'h8793000f ;
			32'h00101560 : data_o = 32'h4398abe7 ;
			32'h00101564 : data_o = 32'h853a43dc ;
			32'h00101568 : data_o = 32'h3f8585be ;
			32'h0010156c : data_o = 32'h000ff797 ;
			32'h00101570 : data_o = 32'haa478793 ;
			32'h00101574 : data_o = 32'h43dc4398 ;
			32'h00101578 : data_o = 32'h45814505 ;
			32'h0010157c : data_o = 32'h00a70633 ;
			32'h00101580 : data_o = 32'h38338832 ;
			32'h00101584 : data_o = 32'h86b300e8 ;
			32'h00101588 : data_o = 32'h07b300b7 ;
			32'h0010158c : data_o = 32'h86be00d8 ;
			32'h00101590 : data_o = 32'h87b68732 ;
			32'h00101594 : data_o = 32'h000ff697 ;
			32'h00101598 : data_o = 32'ha7c68693 ;
			32'h0010159c : data_o = 32'hc2dcc298 ;
			32'h001015a0 : data_o = 32'h40b60001 ;
			32'h001015a4 : data_o = 32'h431642a6 ;
			32'h001015a8 : data_o = 32'h54724386 ;
			32'h001015ac : data_o = 32'h55d25562 ;
			32'h001015b0 : data_o = 32'h56b25642 ;
			32'h001015b4 : data_o = 32'h57925722 ;
			32'h001015b8 : data_o = 32'h48f25802 ;
			32'h001015bc : data_o = 32'h4ed24e62 ;
			32'h001015c0 : data_o = 32'h4fb24f42 ;
			32'h001015c4 : data_o = 32'h00736161 ;
			32'h001015c8 : data_o = 32'h11413020 ;
			32'h001015cc : data_o = 32'h0800c622 ;
			32'h001015d0 : data_o = 32'h44320001 ;
			32'h001015d4 : data_o = 32'h80820141 ;
			32'h001015d8 : data_o = 32'hce221101 ;
			32'h001015dc : data_o = 32'h28371000 ;
			32'h001015e0 : data_o = 32'h08110800 ;
			32'h001015e4 : data_o = 32'h00082803 ;
			32'h001015e8 : data_o = 32'hff042623 ;
			32'h001015ec : data_o = 32'h08002837 ;
			32'h001015f0 : data_o = 32'h00082803 ;
			32'h001015f4 : data_o = 32'hff042423 ;
			32'h001015f8 : data_o = 32'h08002837 ;
			32'h001015fc : data_o = 32'h28030811 ;
			32'h00101600 : data_o = 32'h28830008 ;
			32'h00101604 : data_o = 32'h9ce3fec4 ;
			32'h00101608 : data_o = 32'h2803fd08 ;
			32'h0010160c : data_o = 32'h8542fec4 ;
			32'h00101610 : data_o = 32'h17934581 ;
			32'h00101614 : data_o = 32'h47010005 ;
			32'h00101618 : data_o = 32'hfe842583 ;
			32'h0010161c : data_o = 32'h4681862e ;
			32'h00101620 : data_o = 32'h00c765b3 ;
			32'h00101624 : data_o = 32'hfeb42023 ;
			32'h00101628 : data_o = 32'h22238fd5 ;
			32'h0010162c : data_o = 32'h2703fef4 ;
			32'h00101630 : data_o = 32'h2783fe04 ;
			32'h00101634 : data_o = 32'h853afe44 ;
			32'h00101638 : data_o = 32'h447285be ;
			32'h0010163c : data_o = 32'h80826105 ;
			32'h00101640 : data_o = 32'hc6221141 ;
			32'h00101644 : data_o = 32'hf7970800 ;
			32'h00101648 : data_o = 32'h8793000f ;
			32'h0010164c : data_o = 32'h43989ca7 ;
			32'h00101650 : data_o = 32'h853a43dc ;
			32'h00101654 : data_o = 32'h443285be ;
			32'h00101658 : data_o = 32'h80820141 ;
			32'h0010165c : data_o = 32'hce061101 ;
			32'h00101660 : data_o = 32'h1000cc22 ;
			32'h00101664 : data_o = 32'hfea42423 ;
			32'h00101668 : data_o = 32'hfeb42623 ;
			32'h0010166c : data_o = 32'h000ff797 ;
			32'h00101670 : data_o = 32'h9a478793 ;
			32'h00101674 : data_o = 32'h47014681 ;
			32'h00101678 : data_o = 32'hc3d8c394 ;
			32'h0010167c : data_o = 32'h000ff697 ;
			32'h00101680 : data_o = 32'h99c68693 ;
			32'h00101684 : data_o = 32'hfe842703 ;
			32'h00101688 : data_o = 32'hfec42783 ;
			32'h0010168c : data_o = 32'hc2dcc298 ;
			32'h00101690 : data_o = 32'hfe842503 ;
			32'h00101694 : data_o = 32'hfec42583 ;
			32'h00101698 : data_o = 32'h05133589 ;
			32'h0010169c : data_o = 32'h31e90800 ;
			32'h001016a0 : data_o = 32'h39ed4505 ;
			32'h001016a4 : data_o = 32'h40f20001 ;
			32'h001016a8 : data_o = 32'h61054462 ;
			32'h001016ac : data_o = 32'h11418082 ;
			32'h001016b0 : data_o = 32'h0800c622 ;
			32'h001016b4 : data_o = 32'h08000793 ;
			32'h001016b8 : data_o = 32'h3047b073 ;
			32'h001016bc : data_o = 32'h44320001 ;
			32'h001016c0 : data_o = 32'h80820141 ;
			32'h001016c4 : data_o = 32'hce221101 ;
			32'h001016c8 : data_o = 32'h26231000 ;
			32'h001016cc : data_o = 32'h2423fea4 ;
			32'h001016d0 : data_o = 32'h2783feb4 ;
			32'h001016d4 : data_o = 32'h2703fec4 ;
			32'h001016d8 : data_o = 32'hc398fe84 ;
			32'h001016dc : data_o = 32'h44720001 ;
			32'h001016e0 : data_o = 32'h80826105 ;
			32'h001016e4 : data_o = 32'hce221101 ;
			32'h001016e8 : data_o = 32'h26231000 ;
			32'h001016ec : data_o = 32'h2783fea4 ;
			32'h001016f0 : data_o = 32'h439cfec4 ;
			32'h001016f4 : data_o = 32'h4472853e ;
			32'h001016f8 : data_o = 32'h80826105 ;
			32'h001016fc : data_o = 32'hd6067179 ;
			32'h00101700 : data_o = 32'h1800d422 ;
			32'h00101704 : data_o = 32'hfca42e23 ;
			32'h00101708 : data_o = 32'hfcb42c23 ;
			32'h0010170c : data_o = 32'hfcc42a23 ;
			32'h00101710 : data_o = 32'hfdc42503 ;
			32'h00101714 : data_o = 32'h26233fc1 ;
			32'h00101718 : data_o = 32'h2783fea4 ;
			32'h0010171c : data_o = 32'h4705fd84 ;
			32'h00101720 : data_o = 32'h00f717b3 ;
			32'h00101724 : data_o = 32'hfff7c793 ;
			32'h00101728 : data_o = 32'h2783873e ;
			32'h0010172c : data_o = 32'h8ff9fec4 ;
			32'h00101730 : data_o = 32'hfef42623 ;
			32'h00101734 : data_o = 32'hfd842783 ;
			32'h00101738 : data_o = 32'hfd442703 ;
			32'h0010173c : data_o = 32'h00f717b3 ;
			32'h00101740 : data_o = 32'hfec42703 ;
			32'h00101744 : data_o = 32'h26238fd9 ;
			32'h00101748 : data_o = 32'h2583fef4 ;
			32'h0010174c : data_o = 32'h2503fec4 ;
			32'h00101750 : data_o = 32'h3f8dfdc4 ;
			32'h00101754 : data_o = 32'h50b20001 ;
			32'h00101758 : data_o = 32'h61455422 ;
			32'h0010175c : data_o = 32'h71798082 ;
			32'h00101760 : data_o = 32'hd422d606 ;
			32'h00101764 : data_o = 32'h2e231800 ;
			32'h00101768 : data_o = 32'h2c23fca4 ;
			32'h0010176c : data_o = 32'h2503fcb4 ;
			32'h00101770 : data_o = 32'h3f8dfdc4 ;
			32'h00101774 : data_o = 32'hfea42623 ;
			32'h00101778 : data_o = 32'hfd842783 ;
			32'h0010177c : data_o = 32'hfec42703 ;
			32'h00101780 : data_o = 32'h00f757b3 ;
			32'h00101784 : data_o = 32'h853e8b85 ;
			32'h00101788 : data_o = 32'h542250b2 ;
			32'h0010178c : data_o = 32'h80826145 ;
			32'h00101790 : data_o = 32'hce221101 ;
			32'h00101794 : data_o = 32'h26231000 ;
			32'h00101798 : data_o = 32'h07b7fea4 ;
			32'h0010179c : data_o = 32'h07c17000 ;
			32'h001017a0 : data_o = 32'hfec42703 ;
			32'h001017a4 : data_o = 32'h0001c398 ;
			32'h001017a8 : data_o = 32'h61054472 ;
			32'h001017ac : data_o = 32'h71798082 ;
			32'h001017b0 : data_o = 32'h1800d622 ;
			32'h001017b4 : data_o = 32'hfca42e23 ;
			32'h001017b8 : data_o = 32'hfdc42783 ;
			32'h001017bc : data_o = 32'h0007c783 ;
			32'h001017c0 : data_o = 32'h2783873e ;
			32'h001017c4 : data_o = 32'h0785fdc4 ;
			32'h001017c8 : data_o = 32'h0007c783 ;
			32'h001017cc : data_o = 32'h8f5d07a2 ;
			32'h001017d0 : data_o = 32'hfdc42783 ;
			32'h001017d4 : data_o = 32'hc7830789 ;
			32'h001017d8 : data_o = 32'h07c20007 ;
			32'h001017dc : data_o = 32'h27838f5d ;
			32'h001017e0 : data_o = 32'h078dfdc4 ;
			32'h001017e4 : data_o = 32'h0007c783 ;
			32'h001017e8 : data_o = 32'h8fd907e2 ;
			32'h001017ec : data_o = 32'hfef42623 ;
			32'h001017f0 : data_o = 32'h700007b7 ;
			32'h001017f4 : data_o = 32'h270307e1 ;
			32'h001017f8 : data_o = 32'hc398fec4 ;
			32'h001017fc : data_o = 32'h54320001 ;
			32'h00101800 : data_o = 32'h80826145 ;
			32'h00101804 : data_o = 32'hc6221141 ;
			32'h00101808 : data_o = 32'h07b70800 ;
			32'h0010180c : data_o = 32'h87937000 ;
			32'h00101810 : data_o = 32'h47050207 ;
			32'h00101814 : data_o = 32'h0001c398 ;
			32'h00101818 : data_o = 32'h01414432 ;
			32'h0010181c : data_o = 32'h11418082 ;
			32'h00101820 : data_o = 32'h0800c622 ;
			32'h00101824 : data_o = 32'h07b70001 ;
			32'h00101828 : data_o = 32'h87937000 ;
			32'h0010182c : data_o = 32'h439c0247 ;
			32'h00101830 : data_o = 32'h07b7dbfd ;
			32'h00101834 : data_o = 32'h87937000 ;
			32'h00101838 : data_o = 32'h439c0287 ;
			32'h0010183c : data_o = 32'h4432853e ;
			32'h00101840 : data_o = 32'h80820141 ;
			32'h00101844 : data_o = 32'hc6061141 ;
			32'h00101848 : data_o = 32'h0800c422 ;
			32'h0010184c : data_o = 32'h00020537 ;
			32'h00101850 : data_o = 32'h45053e21 ;
			32'h00101854 : data_o = 32'h07b736a1 ;
			32'h00101858 : data_o = 32'h87937000 ;
			32'h0010185c : data_o = 32'h47050307 ;
			32'h00101860 : data_o = 32'h0001c398 ;
			32'h00101864 : data_o = 32'h442240b2 ;
			32'h00101868 : data_o = 32'h80820141 ;
			32'h0010186c : data_o = 32'hc6061141 ;
			32'h00101870 : data_o = 32'h0800c422 ;
			32'h00101874 : data_o = 32'h700007b7 ;
			32'h00101878 : data_o = 32'h03078793 ;
			32'h0010187c : data_o = 32'h0007a023 ;
			32'h00101880 : data_o = 32'h00020537 ;
			32'h00101884 : data_o = 32'h00013cfd ;
			32'h00101888 : data_o = 32'h442240b2 ;
			32'h0010188c : data_o = 32'h80820141 ;
			32'h00101890 : data_o = 32'hce221101 ;
			32'h00101894 : data_o = 32'h26231000 ;
			32'h00101898 : data_o = 32'h07b7fea4 ;
			32'h0010189c : data_o = 32'h87937000 ;
			32'h001018a0 : data_o = 32'h27030347 ;
			32'h001018a4 : data_o = 32'hc398fec4 ;
			32'h001018a8 : data_o = 32'h44720001 ;
			32'h001018ac : data_o = 32'h80826105 ;
			32'h001018b0 : data_o = 32'hce221101 ;
			32'h001018b4 : data_o = 32'h26231000 ;
			32'h001018b8 : data_o = 32'h07b7fea4 ;
			32'h001018bc : data_o = 32'h87937000 ;
			32'h001018c0 : data_o = 32'h071303c7 ;
			32'h001018c4 : data_o = 32'hc398fec4 ;
			32'h001018c8 : data_o = 32'h44720001 ;
			32'h001018cc : data_o = 32'h80826105 ;
			32'h001018d0 : data_o = 32'hce221101 ;
			32'h001018d4 : data_o = 32'h26231000 ;
			32'h001018d8 : data_o = 32'h07b7fea4 ;
			32'h001018dc : data_o = 32'h87937000 ;
			32'h001018e0 : data_o = 32'h27030387 ;
			32'h001018e4 : data_o = 32'hc398fec4 ;
			32'h001018e8 : data_o = 32'h44720001 ;
			32'h001018ec : data_o = 32'h80826105 ;
			32'h001018f0 : data_o = 32'hc6221141 ;
			32'h001018f4 : data_o = 32'h07b70800 ;
			32'h001018f8 : data_o = 32'h87937000 ;
			32'h001018fc : data_o = 32'h439c0407 ;
			32'h00101900 : data_o = 32'h0ff7f793 ;
			32'h00101904 : data_o = 32'h4432853e ;
			32'h00101908 : data_o = 32'h80820141 ;
			32'h0010190c : data_o = 32'hc6221141 ;
			32'h00101910 : data_o = 32'h07b70800 ;
			32'h00101914 : data_o = 32'h87937000 ;
			32'h00101918 : data_o = 32'h47050447 ;
			32'h0010191c : data_o = 32'h0001c398 ;
			32'h00101920 : data_o = 32'h01414432 ;
			32'h00101924 : data_o = 32'h11418082 ;
			32'h00101928 : data_o = 32'h0800c622 ;
			32'h0010192c : data_o = 32'h700007b7 ;
			32'h00101930 : data_o = 32'h04478793 ;
			32'h00101934 : data_o = 32'h0007a023 ;
			32'h00101938 : data_o = 32'h44320001 ;
			32'h0010193c : data_o = 32'h80820141 ;
			32'h00101940 : data_o = 32'hce221101 ;
			32'h00101944 : data_o = 32'h26231000 ;
			32'h00101948 : data_o = 32'h07b7fea4 ;
			32'h0010194c : data_o = 32'h87937000 ;
			32'h00101950 : data_o = 32'h27030487 ;
			32'h00101954 : data_o = 32'hc398fec4 ;
			32'h00101958 : data_o = 32'h44720001 ;
			32'h0010195c : data_o = 32'h80826105 ;
			32'h00101960 : data_o = 32'hce221101 ;
			32'h00101964 : data_o = 32'h26231000 ;
			32'h00101968 : data_o = 32'h07b7fea4 ;
			32'h0010196c : data_o = 32'h87937000 ;
			32'h00101970 : data_o = 32'h270304c7 ;
			32'h00101974 : data_o = 32'hc398fec4 ;
			32'h00101978 : data_o = 32'h44720001 ;
			32'h0010197c : data_o = 32'h80826105 ;
			32'h00101980 : data_o = 32'hce221101 ;
			32'h00101984 : data_o = 32'h26231000 ;
			32'h00101988 : data_o = 32'h87aefea4 ;
			32'h0010198c : data_o = 32'h05a38732 ;
			32'h00101990 : data_o = 32'h87bafef4 ;
			32'h00101994 : data_o = 32'hfef40523 ;
			32'h00101998 : data_o = 32'hfec42783 ;
			32'h0010199c : data_o = 32'h4703439c ;
			32'h001019a0 : data_o = 32'h0716feb4 ;
			32'h001019a4 : data_o = 32'h06077693 ;
			32'h001019a8 : data_o = 32'h70001737 ;
			32'h001019ac : data_o = 32'h80070713 ;
			32'h001019b0 : data_o = 32'h47038ed9 ;
			32'h001019b4 : data_o = 32'h070afea4 ;
			32'h001019b8 : data_o = 32'h8f558b71 ;
			32'h001019bc : data_o = 32'hfff7c793 ;
			32'h001019c0 : data_o = 32'h0001c31c ;
			32'h001019c4 : data_o = 32'h61054472 ;
			32'h001019c8 : data_o = 32'hf06f8082 ;
			32'h001019cc : data_o = 32'h00939f9f ;
			32'h001019d0 : data_o = 32'h81060000 ;
			32'h001019d4 : data_o = 32'h82068186 ;
			32'h001019d8 : data_o = 32'h83068286 ;
			32'h001019dc : data_o = 32'h84068386 ;
			32'h001019e0 : data_o = 32'h85068486 ;
			32'h001019e4 : data_o = 32'h86068586 ;
			32'h001019e8 : data_o = 32'h87068686 ;
			32'h001019ec : data_o = 32'h88068786 ;
			32'h001019f0 : data_o = 32'h89068886 ;
			32'h001019f4 : data_o = 32'h8a068986 ;
			32'h001019f8 : data_o = 32'h8b068a86 ;
			32'h001019fc : data_o = 32'h8c068b86 ;
			32'h00101a00 : data_o = 32'h8d068c86 ;
			32'h00101a04 : data_o = 32'h8e068d86 ;
			32'h00101a08 : data_o = 32'h8f068e86 ;
			32'h00101a0c : data_o = 32'he1178f86 ;
			32'h00101a10 : data_o = 32'h01130011 ;
			32'h00101a14 : data_o = 32'hed175f21 ;
			32'h00101a18 : data_o = 32'h0d13000f ;
			32'h00101a1c : data_o = 32'hed975f2d ;
			32'h00101a20 : data_o = 32'h8d93000f ;
			32'h00101a24 : data_o = 32'h5763602d ;
			32'h00101a28 : data_o = 32'h202301bd ;
			32'h00101a2c : data_o = 32'h0d11000d ;
			32'h00101a30 : data_o = 32'hffaddde3 ;
			32'h00101a34 : data_o = 32'h45814501 ;
			32'h00101a38 : data_o = 32'hb33fe0ef ;
			32'h00101a3c : data_o = 32'h000202b7 ;
			32'h00101a40 : data_o = 32'h430502a1 ;
			32'h00101a44 : data_o = 32'h0062a023 ;
			32'h00101a48 : data_o = 32'h10500073 ;
			32'h00101a4c : data_o = 32'h47b3bff5 ;
			32'h00101a50 : data_o = 32'h8b8d00b5 ;
			32'h00101a54 : data_o = 32'h00c508b3 ;
			32'h00101a58 : data_o = 32'h478de7b1 ;
			32'h00101a5c : data_o = 32'h04c7f463 ;
			32'h00101a60 : data_o = 32'h00357793 ;
			32'h00101a64 : data_o = 32'hebb9872a ;
			32'h00101a68 : data_o = 32'hffc8f613 ;
			32'h00101a6c : data_o = 32'h40e606b3 ;
			32'h00101a70 : data_o = 32'h02000793 ;
			32'h00101a74 : data_o = 32'h06d7c863 ;
			32'h00101a78 : data_o = 32'h87ba86ae ;
			32'h00101a7c : data_o = 32'h02c77163 ;
			32'h00101a80 : data_o = 32'h0006a803 ;
			32'h00101a84 : data_o = 32'h06910791 ;
			32'h00101a88 : data_o = 32'hff07ae23 ;
			32'h00101a8c : data_o = 32'hfec7eae3 ;
			32'h00101a90 : data_o = 32'hfff60793 ;
			32'h00101a94 : data_o = 32'h9bf18f99 ;
			32'h00101a98 : data_o = 32'h973e0791 ;
			32'h00101a9c : data_o = 32'h666395be ;
			32'h00101aa0 : data_o = 32'h80820117 ;
			32'h00101aa4 : data_o = 32'h7e63872a ;
			32'h00101aa8 : data_o = 32'hc7830315 ;
			32'h00101aac : data_o = 32'h07050005 ;
			32'h00101ab0 : data_o = 32'h0fa30585 ;
			32'h00101ab4 : data_o = 32'h9ae3fef7 ;
			32'h00101ab8 : data_o = 32'h8082fee8 ;
			32'h00101abc : data_o = 32'h0005c683 ;
			32'h00101ac0 : data_o = 32'h77930705 ;
			32'h00101ac4 : data_o = 32'h0fa30037 ;
			32'h00101ac8 : data_o = 32'h0585fed7 ;
			32'h00101acc : data_o = 32'hc683dfd1 ;
			32'h00101ad0 : data_o = 32'h07050005 ;
			32'h00101ad4 : data_o = 32'h00377793 ;
			32'h00101ad8 : data_o = 32'hfed70fa3 ;
			32'h00101adc : data_o = 32'hfff90585 ;
			32'h00101ae0 : data_o = 32'h8082b761 ;
			32'h00101ae4 : data_o = 32'hc6221141 ;
			32'h00101ae8 : data_o = 32'h02000413 ;
			32'h00101aec : data_o = 32'h0005a383 ;
			32'h00101af0 : data_o = 32'h0045a283 ;
			32'h00101af4 : data_o = 32'h0085af83 ;
			32'h00101af8 : data_o = 32'h00c5af03 ;
			32'h00101afc : data_o = 32'h0105ae83 ;
			32'h00101b00 : data_o = 32'h0145ae03 ;
			32'h00101b04 : data_o = 32'h0185a303 ;
			32'h00101b08 : data_o = 32'h01c5a803 ;
			32'h00101b0c : data_o = 32'h07135194 ;
			32'h00101b10 : data_o = 32'h07b30247 ;
			32'h00101b14 : data_o = 32'h2e2340e6 ;
			32'h00101b18 : data_o = 32'h2023fc77 ;
			32'h00101b1c : data_o = 32'h2223fe57 ;
			32'h00101b20 : data_o = 32'h2423fff7 ;
			32'h00101b24 : data_o = 32'h2623ffe7 ;
			32'h00101b28 : data_o = 32'h2823ffd7 ;
			32'h00101b2c : data_o = 32'h2a23ffc7 ;
			32'h00101b30 : data_o = 32'h2c23fe67 ;
			32'h00101b34 : data_o = 32'h2e23ff07 ;
			32'h00101b38 : data_o = 32'h8593fed7 ;
			32'h00101b3c : data_o = 32'h47e30245 ;
			32'h00101b40 : data_o = 32'h86aefaf4 ;
			32'h00101b44 : data_o = 32'h716387ba ;
			32'h00101b48 : data_o = 32'ha80302c7 ;
			32'h00101b4c : data_o = 32'h07910006 ;
			32'h00101b50 : data_o = 32'hae230691 ;
			32'h00101b54 : data_o = 32'heae3ff07 ;
			32'h00101b58 : data_o = 32'h0793fec7 ;
			32'h00101b5c : data_o = 32'h8f99fff6 ;
			32'h00101b60 : data_o = 32'h07919bf1 ;
			32'h00101b64 : data_o = 32'h95be973e ;
			32'h00101b68 : data_o = 32'h01176563 ;
			32'h00101b6c : data_o = 32'h01414432 ;
			32'h00101b70 : data_o = 32'hc7838082 ;
			32'h00101b74 : data_o = 32'h07050005 ;
			32'h00101b78 : data_o = 32'h0fa30585 ;
			32'h00101b7c : data_o = 32'h87e3fef7 ;
			32'h00101b80 : data_o = 32'hc783fee8 ;
			32'h00101b84 : data_o = 32'h07050005 ;
			32'h00101b88 : data_o = 32'h0fa30585 ;
			32'h00101b8c : data_o = 32'h92e3fef7 ;
			32'h00101b90 : data_o = 32'hbfe9fee8 ;
			32'h00101b94 : data_o = 32'h73696854 ;
			32'h00101b98 : data_o = 32'h20736920 ;
			32'h00101b9c : data_o = 32'h20656874 ;
			32'h00101ba0 : data_o = 32'h746f6f62 ;
			32'h00101ba4 : data_o = 32'h64616f6c ;
			32'h00101ba8 : data_o = 32'h0a2e7265 ;
			32'h00101bac : data_o = 32'h00000000 ;
			32'h00101bb0 : data_o = 32'h72617453 ;
			32'h00101bb4 : data_o = 32'h656d2074 ;
			32'h00101bb8 : data_o = 32'h72757361 ;
			32'h00101bbc : data_o = 32'h00000a65 ;
			32'h00101bc0 : data_o = 32'h6d726f46 ;
			32'h00101bc4 : data_o = 32'h20676e69 ;
			32'h00101bc8 : data_o = 32'h62616e45 ;
			32'h00101bcc : data_o = 32'h0a64656c ;
			32'h00101bd0 : data_o = 32'h00000000 ;
			32'h00101bd4 : data_o = 32'h676f7250 ;
			32'h00101bd8 : data_o = 32'h6d6d6172 ;
			32'h00101bdc : data_o = 32'h20676e69 ;
			32'h00101be0 : data_o = 32'h62616e45 ;
			32'h00101be4 : data_o = 32'h0a64656c ;
			32'h00101be8 : data_o = 32'h00000000 ;
			32'h00101bec : data_o = 32'h45534552 ;
			32'h00101bf0 : data_o = 32'h00000a54 ;
			32'h00101bf4 : data_o = 32'h0a544553 ;
			32'h00101bf8 : data_o = 32'h00000000 ;
			32'h00101bfc : data_o = 32'h696e6966 ;
			32'h00101c00 : data_o = 32'h70206873 ;
			32'h00101c04 : data_o = 32'h72676f72 ;
			32'h00101c08 : data_o = 32'h696d6d61 ;
			32'h00101c0c : data_o = 32'h000a676e ;
			32'h00101c10 : data_o = 32'h44414552 ;
			32'h00101c14 : data_o = 32'h0000000a ;
			32'h00101c18 : data_o = 32'h74697277 ;
			32'h00101c1c : data_o = 32'h72652065 ;
			32'h00101c20 : data_o = 32'h73726f72 ;
			32'h00101c24 : data_o = 32'h00203a20 ;
			32'h00101c28 : data_o = 32'h44414552 ;
			32'h00101c2c : data_o = 32'h64647620 ;
			32'h00101c30 : data_o = 32'h00003a20 ;
			32'h00101c34 : data_o = 32'h6f727265 ;
			32'h00101c38 : data_o = 32'h3a207372 ;
			32'h00101c3c : data_o = 32'h00000000 ;
			32'h00101c40 : data_o = 32'h66666964 ;
			32'h00101c44 : data_o = 32'h00003a20 ;
			32'h00101c48 : data_o = 32'h6e696f70 ;
			32'h00101c4c : data_o = 32'h3a207374 ;
			32'h00101c50 : data_o = 32'h00000000 ;
			32'h00101c54 : data_o = 32'h454e4f44 ;
			32'h00101c58 : data_o = 32'h0000000a ;
			32'h00101c5c : data_o = 32'h5e595729 ;
			32'h00101c60 : data_o = 32'h00000000 ;
			32'h00101c64 : data_o = 32'h4f3d2607 ;
			32'h00101c68 : data_o = 32'h7e74695d ;
			32'h00101c6c : data_o = 32'h271b1118 ;
			32'h00101c70 : data_o = 32'h4e453c32 ;
			32'h00101c74 : data_o = 32'h39548bff ;
			32'h00101c78 : data_o = 32'h1b1e232b ;
			32'h00101c7c : data_o = 32'h847f3e7c ;
			32'h00101c80 : data_o = 32'h00000000 ;
			32'h00101c84 : data_o = 32'h63442016 ;
			32'h00101c88 : data_o = 32'hbca9957d ;
			32'h00101c8c : data_o = 32'h664f3209 ;
			32'h00101c90 : data_o = 32'ha4978979 ;
			32'h00101c94 : data_o = 32'hca3e02ff ;
			32'h00101c98 : data_o = 32'hffffffff ;
			32'h00101c9c : data_o = 32'h401eef45 ;
			32'h00101ca0 : data_o = 32'h00000000 ;
			32'h00101ca4 : data_o = 32'h1d181c79 ;
			32'h00101ca8 : data_o = 32'h3c342c25 ;
			32'h00101cac : data_o = 32'h4335240a ;
			32'h00101cb0 : data_o = 32'h665f574e ;
			32'h00101cb4 : data_o = 32'h0c1a5fff ;
			32'h00101cb8 : data_o = 32'h4a342112 ;
			32'h00101cbc : data_o = 32'h2346f5f5 ;
			32'h00101cc0 : data_o = 32'h00000000 ;
			32'h00101cc4 : data_o = 32'h1e21309d ;
			32'h00101cc8 : data_o = 32'h2825221f ;
			32'h00101ccc : data_o = 32'h52391c07 ;
			32'h00101cd0 : data_o = 32'h9d8d7b68 ;
			32'h00101cd4 : data_o = 32'h190655ff ;
			32'h00101cd8 : data_o = 32'hffd28d4d ;
			32'h00101cdc : data_o = 32'h4d524f46 ;
			32'h00101ce0 : data_o = 32'h0000000a ;
			32'h00101ce4 : data_o = 32'h45435845 ;
			32'h00101ce8 : data_o = 32'h4f495450 ;
			32'h00101cec : data_o = 32'h2121214e ;
			32'h00101cf0 : data_o = 32'h0000000a ;
			32'h00101cf4 : data_o = 32'h3d3d3d3d ;
			32'h00101cf8 : data_o = 32'h3d3d3d3d ;
			32'h00101cfc : data_o = 32'h3d3d3d3d ;
			32'h00101d00 : data_o = 32'h0000000a ;
			32'h00101d04 : data_o = 32'h4350454d ;
			32'h00101d08 : data_o = 32'h2020203a ;
			32'h00101d0c : data_o = 32'h00007830 ;
			32'h00101d10 : data_o = 32'h41434d0a ;
			32'h00101d14 : data_o = 32'h3a455355 ;
			32'h00101d18 : data_o = 32'h00783020 ;
			32'h00101d1c : data_o = 32'h56544d0a ;
			32'h00101d20 : data_o = 32'h203a4c41 ;
			32'h00101d24 : data_o = 32'h00783020 ;
			32'h00101d28 : data_o = 32'h00100000 ;
			default : data_o = 32'h00000000 ;
		endcase 
	end
endmodule
