module rom_1p #(
	int Depth, 
 	int DATA_WIDTH = 32, 
 	int ADDR_WIDTH = 32 
 ) (
	input logic clk_i, 
	input logic req_i, 
	input logic [ADDR_WIDTH-1:0] addr_i, 
	output logic [DATA_WIDTH-1:0] data_o 
 );
	always_ff @(posedge clk_i) begin
		case (addr_i)
			32'h00100000 : data_o = 32'h25a0006f ;
			32'h00100004 : data_o = 32'h2560006f ;
			32'h00100008 : data_o = 32'h2520006f ;
			32'h0010000c : data_o = 32'h24e0006f ;
			32'h00100010 : data_o = 32'h24a0006f ;
			32'h00100014 : data_o = 32'h2460006f ;
			32'h00100018 : data_o = 32'h2420006f ;
			32'h0010001c : data_o = 32'h23e0006f ;
			32'h00100020 : data_o = 32'h23a0006f ;
			32'h00100024 : data_o = 32'h2360006f ;
			32'h00100028 : data_o = 32'h2320006f ;
			32'h0010002c : data_o = 32'h22e0006f ;
			32'h00100030 : data_o = 32'h22a0006f ;
			32'h00100034 : data_o = 32'h2260006f ;
			32'h00100038 : data_o = 32'h2220006f ;
			32'h0010003c : data_o = 32'h21e0006f ;
			32'h00100040 : data_o = 32'h21a0006f ;
			32'h00100044 : data_o = 32'h0400006f ;
			32'h00100048 : data_o = 32'h2120006f ;
			32'h0010004c : data_o = 32'h20e0006f ;
			32'h00100050 : data_o = 32'h20a0006f ;
			32'h00100054 : data_o = 32'h2060006f ;
			32'h00100058 : data_o = 32'h2020006f ;
			32'h0010005c : data_o = 32'h1fe0006f ;
			32'h00100060 : data_o = 32'h1fa0006f ;
			32'h00100064 : data_o = 32'h1f60006f ;
			32'h00100068 : data_o = 32'h1f20006f ;
			32'h0010006c : data_o = 32'h1ee0006f ;
			32'h00100070 : data_o = 32'h1ea0006f ;
			32'h00100074 : data_o = 32'h1e60006f ;
			32'h00100078 : data_o = 32'h1e20006f ;
			32'h0010007c : data_o = 32'h1de0006f ;
			32'h00100080 : data_o = 32'h46c0006f ;
			32'h00100084 : data_o = 32'hde067139 ;
			32'h00100088 : data_o = 32'hda1adc16 ;
			32'h0010008c : data_o = 32'hd62ad81e ;
			32'h00100090 : data_o = 32'hd232d42e ;
			32'h00100094 : data_o = 32'hce3ad036 ;
			32'h00100098 : data_o = 32'hca42cc3e ;
			32'h0010009c : data_o = 32'hc672c846 ;
			32'h001000a0 : data_o = 32'hc27ac476 ;
			32'h001000a4 : data_o = 32'h2e51c07e ;
			32'h001000a8 : data_o = 32'h00100797 ;
			32'h001000ac : data_o = 32'hf6a7a623 ;
			32'h001000b0 : data_o = 32'h07174785 ;
			32'h001000b4 : data_o = 32'h2f230010 ;
			32'h001000b8 : data_o = 32'h50f2f4f7 ;
			32'h001000bc : data_o = 32'h535252e2 ;
			32'h001000c0 : data_o = 32'h553253c2 ;
			32'h001000c4 : data_o = 32'h561255a2 ;
			32'h001000c8 : data_o = 32'h47725682 ;
			32'h001000cc : data_o = 32'h485247e2 ;
			32'h001000d0 : data_o = 32'h4e3248c2 ;
			32'h001000d4 : data_o = 32'h4f124ea2 ;
			32'h001000d8 : data_o = 32'h61214f82 ;
			32'h001000dc : data_o = 32'h30200073 ;
			32'h001000e0 : data_o = 32'hc6061141 ;
			32'h001000e4 : data_o = 32'h08000737 ;
			32'h001000e8 : data_o = 32'haaaab7b7 ;
			32'h001000ec : data_o = 32'haaa78793 ;
			32'h001000f0 : data_o = 32'h0517c31c ;
			32'h001000f4 : data_o = 32'h05130000 ;
			32'h001000f8 : data_o = 32'h208548e5 ;
			32'h001000fc : data_o = 32'h00000517 ;
			32'h00100100 : data_o = 32'h4a450513 ;
			32'h00100104 : data_o = 32'h20912899 ;
			32'h00100108 : data_o = 32'h0ff57513 ;
			32'h0010010c : data_o = 32'h05172811 ;
			32'h00100110 : data_o = 32'h05130000 ;
			32'h00100114 : data_o = 32'h209149a5 ;
			32'h00100118 : data_o = 32'h40b24501 ;
			32'h0010011c : data_o = 32'h80820141 ;
			32'h00100120 : data_o = 32'hc6061141 ;
			32'h00100124 : data_o = 32'h842ac422 ;
			32'h00100128 : data_o = 32'h0b6347a9 ;
			32'h0010012c : data_o = 32'h85a200f5 ;
			32'h00100130 : data_o = 32'h80001537 ;
			32'h00100134 : data_o = 32'h85222a51 ;
			32'h00100138 : data_o = 32'h442240b2 ;
			32'h0010013c : data_o = 32'h80820141 ;
			32'h00100140 : data_o = 32'h153745b5 ;
			32'h00100144 : data_o = 32'h22498000 ;
			32'h00100148 : data_o = 32'h1141b7dd ;
			32'h0010014c : data_o = 32'h1537c606 ;
			32'h00100150 : data_o = 32'h22a58000 ;
			32'h00100154 : data_o = 32'h014140b2 ;
			32'h00100158 : data_o = 32'h11418082 ;
			32'h0010015c : data_o = 32'hc422c606 ;
			32'h00100160 : data_o = 32'h4503842a ;
			32'h00100164 : data_o = 32'hc5110005 ;
			32'h00100168 : data_o = 32'h3f5d0405 ;
			32'h0010016c : data_o = 32'h00044503 ;
			32'h00100170 : data_o = 32'h4501fd65 ;
			32'h00100174 : data_o = 32'h442240b2 ;
			32'h00100178 : data_o = 32'h80820141 ;
			32'h0010017c : data_o = 32'hc6061141 ;
			32'h00100180 : data_o = 32'hc226c422 ;
			32'h00100184 : data_o = 32'h842ac04a ;
			32'h00100188 : data_o = 32'h492544a1 ;
			32'h0010018c : data_o = 32'h0513a039 ;
			32'h00100190 : data_o = 32'h37790375 ;
			32'h00100194 : data_o = 32'h14fd0412 ;
			32'h00100198 : data_o = 32'h5513c889 ;
			32'h0010019c : data_o = 32'h48e301c4 ;
			32'h001001a0 : data_o = 32'h0513fea9 ;
			32'h001001a4 : data_o = 32'h3fad0305 ;
			32'h001001a8 : data_o = 32'h40b2b7f5 ;
			32'h001001ac : data_o = 32'h44924422 ;
			32'h001001b0 : data_o = 32'h01414902 ;
			32'h001001b4 : data_o = 32'h07b78082 ;
			32'h001001b8 : data_o = 32'h47050002 ;
			32'h001001bc : data_o = 32'h8082c798 ;
			32'h001001c0 : data_o = 32'h34102573 ;
			32'h001001c4 : data_o = 32'h25738082 ;
			32'h001001c8 : data_o = 32'h80823420 ;
			32'h001001cc : data_o = 32'h34302573 ;
			32'h001001d0 : data_o = 32'h25738082 ;
			32'h001001d4 : data_o = 32'h8082b000 ;
			32'h001001d8 : data_o = 32'hb0001073 ;
			32'h001001dc : data_o = 32'h47fd8082 ;
			32'h001001e0 : data_o = 32'h04a7ec63 ;
			32'h001001e4 : data_o = 32'h0717050a ;
			32'h001001e8 : data_o = 32'h27030010 ;
			32'h001001ec : data_o = 32'h972ae1a7 ;
			32'h001001f0 : data_o = 32'h07b78d99 ;
			32'h001001f4 : data_o = 32'h97ae0008 ;
			32'h001001f8 : data_o = 32'h001006b7 ;
			32'h001001fc : data_o = 32'hfe634509 ;
			32'h00100200 : data_o = 32'h979302d7 ;
			32'h00100204 : data_o = 32'h06b70145 ;
			32'h00100208 : data_o = 32'h8ff57fe0 ;
			32'h0010020c : data_o = 32'h00b59693 ;
			32'h00100210 : data_o = 32'h80000637 ;
			32'h00100214 : data_o = 32'h8fd58ef1 ;
			32'h00100218 : data_o = 32'h000ff6b7 ;
			32'h0010021c : data_o = 32'h8fd58eed ;
			32'h00100220 : data_o = 32'h06b705a6 ;
			32'h00100224 : data_o = 32'h8df50010 ;
			32'h00100228 : data_o = 32'he7938fcd ;
			32'h0010022c : data_o = 32'hc31c06f7 ;
			32'h00100230 : data_o = 32'h0000100f ;
			32'h00100234 : data_o = 32'h80824501 ;
			32'h00100238 : data_o = 32'h80824505 ;
			32'h0010023c : data_o = 32'h30452073 ;
			32'h00100240 : data_o = 32'h30738082 ;
			32'h00100244 : data_o = 32'h80823045 ;
			32'h00100248 : data_o = 32'h47a1c509 ;
			32'h0010024c : data_o = 32'h3007a073 ;
			32'h00100250 : data_o = 32'h47a18082 ;
			32'h00100254 : data_o = 32'h3007b073 ;
			32'h00100258 : data_o = 32'h11418082 ;
			32'h0010025c : data_o = 32'h0517c606 ;
			32'h00100260 : data_o = 32'h05130000 ;
			32'h00100264 : data_o = 32'h3dd535e5 ;
			32'h00100268 : data_o = 32'h00000517 ;
			32'h0010026c : data_o = 32'h36450513 ;
			32'h00100270 : data_o = 32'h051735ed ;
			32'h00100274 : data_o = 32'h05130000 ;
			32'h00100278 : data_o = 32'h35c536a5 ;
			32'h0010027c : data_o = 32'h34102573 ;
			32'h00100280 : data_o = 32'h05173df5 ;
			32'h00100284 : data_o = 32'h05130000 ;
			32'h00100288 : data_o = 32'h3dc13665 ;
			32'h0010028c : data_o = 32'h34202573 ;
			32'h00100290 : data_o = 32'h051735f5 ;
			32'h00100294 : data_o = 32'h05130000 ;
			32'h00100298 : data_o = 32'h35c13625 ;
			32'h0010029c : data_o = 32'h34302573 ;
			32'h001002a0 : data_o = 32'h45293df1 ;
			32'h001002a4 : data_o = 32'ha0013db5 ;
			32'h001002a8 : data_o = 32'hc6061141 ;
			32'h001002ac : data_o = 32'h37796541 ;
			32'h001002b0 : data_o = 32'h3f594505 ;
			32'h001002b4 : data_o = 32'h014140b2 ;
			32'h001002b8 : data_o = 32'h451c8082 ;
			32'h001002bc : data_o = 32'he3998b85 ;
			32'h001002c0 : data_o = 32'h80824108 ;
			32'h001002c4 : data_o = 32'h8082557d ;
			32'h001002c8 : data_o = 32'h8b89451c ;
			32'h001002cc : data_o = 32'hc14cfff5 ;
			32'h001002d0 : data_o = 32'h27b78082 ;
			32'h001002d4 : data_o = 32'h577d0800 ;
			32'h001002d8 : data_o = 32'hc7ccc798 ;
			32'h001002dc : data_o = 32'h8082c788 ;
			32'h001002e0 : data_o = 32'h27b78082 ;
			32'h001002e4 : data_o = 32'h43cc0800 ;
			32'h001002e8 : data_o = 32'h43d84388 ;
			32'h001002ec : data_o = 32'hfeb71de3 ;
			32'h001002f0 : data_o = 32'h715d8082 ;
			32'h001002f4 : data_o = 32'hc496c686 ;
			32'h001002f8 : data_o = 32'hc09ec29a ;
			32'h001002fc : data_o = 32'hdc26de22 ;
			32'h00100300 : data_o = 32'hd82eda2a ;
			32'h00100304 : data_o = 32'hd436d632 ;
			32'h00100308 : data_o = 32'hd03ed23a ;
			32'h0010030c : data_o = 32'hcc46ce42 ;
			32'h00100310 : data_o = 32'hc876ca72 ;
			32'h00100314 : data_o = 32'hc47ec67a ;
			32'h00100318 : data_o = 32'h00100797 ;
			32'h0010031c : data_o = 32'hd0078793 ;
			32'h00100320 : data_o = 32'h43c44380 ;
			32'h00100324 : data_o = 32'h95223f7d ;
			32'h00100328 : data_o = 32'h00853433 ;
			32'h0010032c : data_o = 32'h95a295a6 ;
			32'h00100330 : data_o = 32'h0597374d ;
			32'h00100334 : data_o = 32'h85930010 ;
			32'h00100338 : data_o = 32'h4180cee5 ;
			32'h0010033c : data_o = 32'h051341c4 ;
			32'h00100340 : data_o = 32'h36330014 ;
			32'h00100344 : data_o = 32'h07b30085 ;
			32'h00100348 : data_o = 32'hc1880096 ;
			32'h0010034c : data_o = 32'h40b6c1dc ;
			32'h00100350 : data_o = 32'h431642a6 ;
			32'h00100354 : data_o = 32'h54724386 ;
			32'h00100358 : data_o = 32'h555254e2 ;
			32'h0010035c : data_o = 32'h563255c2 ;
			32'h00100360 : data_o = 32'h571256a2 ;
			32'h00100364 : data_o = 32'h48725782 ;
			32'h00100368 : data_o = 32'h4e5248e2 ;
			32'h0010036c : data_o = 32'h4f324ec2 ;
			32'h00100370 : data_o = 32'h61614fa2 ;
			32'h00100374 : data_o = 32'h30200073 ;
			32'h00100378 : data_o = 32'h00100797 ;
			32'h0010037c : data_o = 32'hca878793 ;
			32'h00100380 : data_o = 32'h43cc4388 ;
			32'h00100384 : data_o = 32'h11418082 ;
			32'h00100388 : data_o = 32'hc422c606 ;
			32'h0010038c : data_o = 32'h842ac226 ;
			32'h00100390 : data_o = 32'h079784ae ;
			32'h00100394 : data_o = 32'h87930010 ;
			32'h00100398 : data_o = 32'h4681c8e7 ;
			32'h0010039c : data_o = 32'hc3944701 ;
			32'h001003a0 : data_o = 32'h0797c3d8 ;
			32'h001003a4 : data_o = 32'h87930010 ;
			32'h001003a8 : data_o = 32'hc388c767 ;
			32'h001003ac : data_o = 32'h3f15c3cc ;
			32'h001003b0 : data_o = 32'h34339522 ;
			32'h001003b4 : data_o = 32'h95a60085 ;
			32'h001003b8 : data_o = 32'h3f2195a2 ;
			32'h001003bc : data_o = 32'h08000513 ;
			32'h001003c0 : data_o = 32'h45053db5 ;
			32'h001003c4 : data_o = 32'h40b23551 ;
			32'h001003c8 : data_o = 32'h44924422 ;
			32'h001003cc : data_o = 32'h80820141 ;
			32'h001003d0 : data_o = 32'h08000793 ;
			32'h001003d4 : data_o = 32'h3047b073 ;
			32'h001003d8 : data_o = 32'hc10c8082 ;
			32'h001003dc : data_o = 32'h41088082 ;
			32'h001003e0 : data_o = 32'h41188082 ;
			32'h001003e4 : data_o = 32'h97b34785 ;
			32'h001003e8 : data_o = 32'hc79300b7 ;
			32'h001003ec : data_o = 32'h8ff9fff7 ;
			32'h001003f0 : data_o = 32'h00b61633 ;
			32'h001003f4 : data_o = 32'hc1108e5d ;
			32'h001003f8 : data_o = 32'h41088082 ;
			32'h001003fc : data_o = 32'h00b55533 ;
			32'h00100400 : data_o = 32'h80828905 ;
			32'h00100404 : data_o = 32'h700007b7 ;
			32'h00100408 : data_o = 32'h8082cb88 ;
			32'h0010040c : data_o = 32'h00154783 ;
			32'h00100410 : data_o = 32'h470307a2 ;
			32'h00100414 : data_o = 32'h07420025 ;
			32'h00100418 : data_o = 32'h47038fd9 ;
			32'h0010041c : data_o = 32'h8fd90005 ;
			32'h00100420 : data_o = 32'h00354703 ;
			32'h00100424 : data_o = 32'h8fd90762 ;
			32'h00100428 : data_o = 32'h70000737 ;
			32'h0010042c : data_o = 32'h8082cf1c ;
			32'h00100430 : data_o = 32'h700007b7 ;
			32'h00100434 : data_o = 32'hd3984705 ;
			32'h00100438 : data_o = 32'h07378082 ;
			32'h0010043c : data_o = 32'h535c7000 ;
			32'h00100440 : data_o = 32'h07b7dffd ;
			32'h00100444 : data_o = 32'h57887000 ;
			32'h00100448 : data_o = 32'h11418082 ;
			32'h0010044c : data_o = 32'h0537c606 ;
			32'h00100450 : data_o = 32'h33ed0002 ;
			32'h00100454 : data_o = 32'h3bcd4505 ;
			32'h00100458 : data_o = 32'h700007b7 ;
			32'h0010045c : data_o = 32'hdb984705 ;
			32'h00100460 : data_o = 32'h014140b2 ;
			32'h00100464 : data_o = 32'h11418082 ;
			32'h00100468 : data_o = 32'h07b7c606 ;
			32'h0010046c : data_o = 32'ha8237000 ;
			32'h00100470 : data_o = 32'h05370207 ;
			32'h00100474 : data_o = 32'h33f10002 ;
			32'h00100478 : data_o = 32'h014140b2 ;
			32'h0010047c : data_o = 32'h07b78082 ;
			32'h00100480 : data_o = 32'hdbc87000 ;
			32'h00100484 : data_o = 32'h11418082 ;
			32'h00100488 : data_o = 32'h07b70078 ;
			32'h0010048c : data_o = 32'hdfd87000 ;
			32'h00100490 : data_o = 32'h80820141 ;
			32'h00100494 : data_o = 32'h700007b7 ;
			32'h00100498 : data_o = 32'h8082df88 ;
			32'h0010049c : data_o = 32'h700007b7 ;
			32'h001004a0 : data_o = 32'h751343a8 ;
			32'h001004a4 : data_o = 32'h80820ff5 ;
			32'h001004a8 : data_o = 32'h700007b7 ;
			32'h001004ac : data_o = 32'hc3f84705 ;
			32'h001004b0 : data_o = 32'h07b78082 ;
			32'h001004b4 : data_o = 32'ha2237000 ;
			32'h001004b8 : data_o = 32'h80820407 ;
			32'h001004bc : data_o = 32'h700007b7 ;
			32'h001004c0 : data_o = 32'h8082c7a8 ;
			32'h001004c4 : data_o = 32'h700007b7 ;
			32'h001004c8 : data_o = 32'h8082c7e8 ;
			32'h001004cc : data_o = 32'h89e1058e ;
			32'h001004d0 : data_o = 32'h8dd18a15 ;
			32'h001004d4 : data_o = 32'h700017b7 ;
			32'h001004d8 : data_o = 32'h80078793 ;
			32'h001004dc : data_o = 32'h411c8ddd ;
			32'h001004e0 : data_o = 32'hfff7c793 ;
			32'h001004e4 : data_o = 32'h8082c19c ;
			32'h001004e8 : data_o = 32'hd73ff06f ;
			32'h001004ec : data_o = 32'h00000093 ;
			32'h001004f0 : data_o = 32'h81868106 ;
			32'h001004f4 : data_o = 32'h82868206 ;
			32'h001004f8 : data_o = 32'h83868306 ;
			32'h001004fc : data_o = 32'h84868406 ;
			32'h00100500 : data_o = 32'h85868506 ;
			32'h00100504 : data_o = 32'h86868606 ;
			32'h00100508 : data_o = 32'h87868706 ;
			32'h0010050c : data_o = 32'h88868806 ;
			32'h00100510 : data_o = 32'h89868906 ;
			32'h00100514 : data_o = 32'h8a868a06 ;
			32'h00100518 : data_o = 32'h8b868b06 ;
			32'h0010051c : data_o = 32'h8c868c06 ;
			32'h00100520 : data_o = 32'h8d868d06 ;
			32'h00100524 : data_o = 32'h8e868e06 ;
			32'h00100528 : data_o = 32'h8f868f06 ;
			32'h0010052c : data_o = 32'h00110117 ;
			32'h00100530 : data_o = 32'had410113 ;
			32'h00100534 : data_o = 32'h00100d17 ;
			32'h00100538 : data_o = 32'had4d0d13 ;
			32'h0010053c : data_o = 32'h00100d97 ;
			32'h00100540 : data_o = 32'haecd8d93 ;
			32'h00100544 : data_o = 32'h01bd5763 ;
			32'h00100548 : data_o = 32'h000d2023 ;
			32'h0010054c : data_o = 32'hdde30d11 ;
			32'h00100550 : data_o = 32'h4501ffad ;
			32'h00100554 : data_o = 32'hf0ef4581 ;
			32'h00100558 : data_o = 32'h02b7b8bf ;
			32'h0010055c : data_o = 32'h02a10002 ;
			32'h00100560 : data_o = 32'ha0234305 ;
			32'h00100564 : data_o = 32'h00730062 ;
			32'h00100568 : data_o = 32'hbff51050 ;
			32'h0010056c : data_o = 32'h00455845 ;
			32'h00100570 : data_o = 32'h5a495300 ;
			32'h00100574 : data_o = 32'h48430045 ;
			32'h00100578 : data_o = 32'h4600534b ;
			32'h0010057c : data_o = 32'h0048534c ;
			32'h00100580 : data_o = 32'h200a0a0a ;
			32'h00100584 : data_o = 32'h414e4950 ;
			32'h00100588 : data_o = 32'h4c505049 ;
			32'h0010058c : data_o = 32'h4f422045 ;
			32'h00100590 : data_o = 32'h4f4c544f ;
			32'h00100594 : data_o = 32'h52454441 ;
			32'h00100598 : data_o = 32'h0a0a0a20 ;
			32'h0010059c : data_o = 32'h00000000 ;
			32'h001005a0 : data_o = 32'h444d430a ;
			32'h001005a4 : data_o = 32'h00203e3a ;
			32'h001005a8 : data_o = 32'h20646d63 ;
			32'h001005ac : data_o = 32'h6c6c6577 ;
			32'h001005b0 : data_o = 32'h63657220 ;
			32'h001005b4 : data_o = 32'h65766965 ;
			32'h001005b8 : data_o = 32'h00000a64 ;
			32'h001005bc : data_o = 32'h45435845 ;
			32'h001005c0 : data_o = 32'h4f495450 ;
			32'h001005c4 : data_o = 32'h2121214e ;
			32'h001005c8 : data_o = 32'h0000000a ;
			32'h001005cc : data_o = 32'h3d3d3d3d ;
			32'h001005d0 : data_o = 32'h3d3d3d3d ;
			32'h001005d4 : data_o = 32'h3d3d3d3d ;
			32'h001005d8 : data_o = 32'h0000000a ;
			32'h001005dc : data_o = 32'h4350454d ;
			32'h001005e0 : data_o = 32'h2020203a ;
			32'h001005e4 : data_o = 32'h00007830 ;
			32'h001005e8 : data_o = 32'h41434d0a ;
			32'h001005ec : data_o = 32'h3a455355 ;
			32'h001005f0 : data_o = 32'h00783020 ;
			32'h001005f4 : data_o = 32'h56544d0a ;
			32'h001005f8 : data_o = 32'h203a4c41 ;
			32'h001005fc : data_o = 32'h00783020 ;
			32'h00100600 : data_o = 32'h00100000 ;
			default : data_o = 32'h00000000 ;
		endcase 
	end
endmodule
