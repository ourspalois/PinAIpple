module rom_1p #(
	int Depth, 
 	int DATA_WIDTH = 32, 
 	int ADDR_WIDTH = 32 
 ) (
	input logic clk_i, 
	input logic req_i, 
	input logic [ADDR_WIDTH-1:0] addr_i, 
	output logic [DATA_WIDTH-1:0] data_o 
 );
	always_ff @(posedge clk_i) begin
		case (addr_i)
			32'h00100000 : data_o = 32'h6440006f ;
			32'h00100004 : data_o = 32'h6400006f ;
			32'h00100008 : data_o = 32'h63c0006f ;
			32'h0010000c : data_o = 32'h6380006f ;
			32'h00100010 : data_o = 32'h6340006f ;
			32'h00100014 : data_o = 32'h6300006f ;
			32'h00100018 : data_o = 32'h62c0006f ;
			32'h0010001c : data_o = 32'h6280006f ;
			32'h00100020 : data_o = 32'h6240006f ;
			32'h00100024 : data_o = 32'h6200006f ;
			32'h00100028 : data_o = 32'h61c0006f ;
			32'h0010002c : data_o = 32'h6180006f ;
			32'h00100030 : data_o = 32'h6140006f ;
			32'h00100034 : data_o = 32'h6100006f ;
			32'h00100038 : data_o = 32'h60c0006f ;
			32'h0010003c : data_o = 32'h6080006f ;
			32'h00100040 : data_o = 32'h6040006f ;
			32'h00100044 : data_o = 32'h0400006f ;
			32'h00100048 : data_o = 32'h5fc0006f ;
			32'h0010004c : data_o = 32'h5f80006f ;
			32'h00100050 : data_o = 32'h5f40006f ;
			32'h00100054 : data_o = 32'h5f00006f ;
			32'h00100058 : data_o = 32'h5ec0006f ;
			32'h0010005c : data_o = 32'h5e80006f ;
			32'h00100060 : data_o = 32'h5e40006f ;
			32'h00100064 : data_o = 32'h5e00006f ;
			32'h00100068 : data_o = 32'h5dc0006f ;
			32'h0010006c : data_o = 32'h5d80006f ;
			32'h00100070 : data_o = 32'h5d40006f ;
			32'h00100074 : data_o = 32'h5d00006f ;
			32'h00100078 : data_o = 32'h5cc0006f ;
			32'h0010007c : data_o = 32'h5c80006f ;
			32'h00100080 : data_o = 32'h3cf0006f ;
			32'h00100084 : data_o = 32'hc686715d ;
			32'h00100088 : data_o = 32'hc29ac496 ;
			32'h0010008c : data_o = 32'hde22c09e ;
			32'h00100090 : data_o = 32'hda2edc2a ;
			32'h00100094 : data_o = 32'hd636d832 ;
			32'h00100098 : data_o = 32'hd23ed43a ;
			32'h0010009c : data_o = 32'hce46d042 ;
			32'h001000a0 : data_o = 32'hca76cc72 ;
			32'h001000a4 : data_o = 32'hc67ec87a ;
			32'h001000a8 : data_o = 32'h00ef0880 ;
			32'h001000ac : data_o = 32'h872a1f70 ;
			32'h001000b0 : data_o = 32'h00100797 ;
			32'h001000b4 : data_o = 32'hf5878793 ;
			32'h001000b8 : data_o = 32'h0797c398 ;
			32'h001000bc : data_o = 32'h87930010 ;
			32'h001000c0 : data_o = 32'h4705f527 ;
			32'h001000c4 : data_o = 32'h0001c398 ;
			32'h001000c8 : data_o = 32'h42a640b6 ;
			32'h001000cc : data_o = 32'h43864316 ;
			32'h001000d0 : data_o = 32'h55625472 ;
			32'h001000d4 : data_o = 32'h564255d2 ;
			32'h001000d8 : data_o = 32'h572256b2 ;
			32'h001000dc : data_o = 32'h58025792 ;
			32'h001000e0 : data_o = 32'h4e6248f2 ;
			32'h001000e4 : data_o = 32'h4f424ed2 ;
			32'h001000e8 : data_o = 32'h61614fb2 ;
			32'h001000ec : data_o = 32'h30200073 ;
			32'h001000f0 : data_o = 32'hc6061141 ;
			32'h001000f4 : data_o = 32'h0800c422 ;
			32'h001000f8 : data_o = 32'h800007b7 ;
			32'h001000fc : data_o = 32'hc3984705 ;
			32'h00100100 : data_o = 32'h07400513 ;
			32'h00100104 : data_o = 32'h05132479 ;
			32'h00100108 : data_o = 32'h24610650 ;
			32'h0010010c : data_o = 32'h07300513 ;
			32'h00100110 : data_o = 32'h05132449 ;
			32'h00100114 : data_o = 32'h2cb50740 ;
			32'h00100118 : data_o = 32'h2ca54529 ;
			32'h0010011c : data_o = 32'h0000100f ;
			32'h00100120 : data_o = 32'h22094501 ;
			32'h00100124 : data_o = 32'h28fd4505 ;
			32'h00100128 : data_o = 32'h28ed4509 ;
			32'h0010012c : data_o = 32'h28dd450d ;
			32'h00100130 : data_o = 32'h0000100f ;
			32'h00100134 : data_o = 32'h06500513 ;
			32'h00100138 : data_o = 32'h05132ca9 ;
			32'h0010013c : data_o = 32'h2c9106e0 ;
			32'h00100140 : data_o = 32'h06400513 ;
			32'h00100144 : data_o = 32'h452924b9 ;
			32'h00100148 : data_o = 32'h07b724a9 ;
			32'h0010014c : data_o = 32'h47098000 ;
			32'h00100150 : data_o = 32'h4781c398 ;
			32'h00100154 : data_o = 32'h40b2853e ;
			32'h00100158 : data_o = 32'h01414422 ;
			32'h0010015c : data_o = 32'h71798082 ;
			32'h00100160 : data_o = 32'h1800d622 ;
			32'h00100164 : data_o = 32'hfca42e23 ;
			32'h00100168 : data_o = 32'hfcb42c23 ;
			32'h0010016c : data_o = 32'hfe042623 ;
			32'h00100170 : data_o = 32'h2783a089 ;
			32'h00100174 : data_o = 32'h2703fec4 ;
			32'h00100178 : data_o = 32'h57b3fdc4 ;
			32'h0010017c : data_o = 32'h8b8500f7 ;
			32'h00100180 : data_o = 32'h2783cb99 ;
			32'h00100184 : data_o = 32'h2703fec4 ;
			32'h00100188 : data_o = 32'h97bafd84 ;
			32'h0010018c : data_o = 32'h03100713 ;
			32'h00100190 : data_o = 32'h00e78023 ;
			32'h00100194 : data_o = 32'h2783a811 ;
			32'h00100198 : data_o = 32'h2703fec4 ;
			32'h0010019c : data_o = 32'h97bafd84 ;
			32'h001001a0 : data_o = 32'h03000713 ;
			32'h001001a4 : data_o = 32'h00e78023 ;
			32'h001001a8 : data_o = 32'hfec42783 ;
			32'h001001ac : data_o = 32'h26230785 ;
			32'h001001b0 : data_o = 32'h2703fef4 ;
			32'h001001b4 : data_o = 32'h47fdfec4 ;
			32'h001001b8 : data_o = 32'hfae7dde3 ;
			32'h001001bc : data_o = 32'hfd842783 ;
			32'h001001c0 : data_o = 32'h02078793 ;
			32'h001001c4 : data_o = 32'h00078023 ;
			32'h001001c8 : data_o = 32'h54320001 ;
			32'h001001cc : data_o = 32'h80826145 ;
			32'h001001d0 : data_o = 32'hce221101 ;
			32'h001001d4 : data_o = 32'h26231000 ;
			32'h001001d8 : data_o = 32'h2703fea4 ;
			32'h001001dc : data_o = 32'h07b7fec4 ;
			32'h001001e0 : data_o = 32'h87931c00 ;
			32'h001001e4 : data_o = 32'h97ba2007 ;
			32'h001001e8 : data_o = 32'h439c078a ;
			32'h001001ec : data_o = 32'h4472853e ;
			32'h001001f0 : data_o = 32'h80826105 ;
			32'h001001f4 : data_o = 32'hce221101 ;
			32'h001001f8 : data_o = 32'h26231000 ;
			32'h001001fc : data_o = 32'h2423fea4 ;
			32'h00100200 : data_o = 32'h2783feb4 ;
			32'h00100204 : data_o = 32'h2703fe84 ;
			32'h00100208 : data_o = 32'h57b3fec4 ;
			32'h0010020c : data_o = 32'h8b8500f7 ;
			32'h00100210 : data_o = 32'h0793c781 ;
			32'h00100214 : data_o = 32'ha0190310 ;
			32'h00100218 : data_o = 32'h03000793 ;
			32'h0010021c : data_o = 32'h4472853e ;
			32'h00100220 : data_o = 32'h80826105 ;
			32'h00100224 : data_o = 32'hc686715d ;
			32'h00100228 : data_o = 32'hc2a6c4a2 ;
			32'h0010022c : data_o = 32'h2e230880 ;
			32'h00100230 : data_o = 32'h2703faa4 ;
			32'h00100234 : data_o = 32'h478dfbc4 ;
			32'h00100238 : data_o = 32'h00e7f463 ;
			32'h0010023c : data_o = 32'ha2a10001 ;
			32'h00100240 : data_o = 32'hfe042623 ;
			32'h00100244 : data_o = 32'h2783a0a5 ;
			32'h00100248 : data_o = 32'h9713fec4 ;
			32'h0010024c : data_o = 32'h27830027 ;
			32'h00100250 : data_o = 32'h97bafbc4 ;
			32'h00100254 : data_o = 32'h00179713 ;
			32'h00100258 : data_o = 32'hfec42783 ;
			32'h0010025c : data_o = 32'h00179493 ;
			32'h00100260 : data_o = 32'h37bd853a ;
			32'h00100264 : data_o = 32'h9793872a ;
			32'h00100268 : data_o = 32'h17c10024 ;
			32'h0010026c : data_o = 32'ha82397a2 ;
			32'h00100270 : data_o = 32'h2783fce7 ;
			32'h00100274 : data_o = 32'h9713fec4 ;
			32'h00100278 : data_o = 32'h27830027 ;
			32'h0010027c : data_o = 32'h97bafbc4 ;
			32'h00100280 : data_o = 32'h87130786 ;
			32'h00100284 : data_o = 32'h27830017 ;
			32'h00100288 : data_o = 32'h0786fec4 ;
			32'h0010028c : data_o = 32'h00178493 ;
			32'h00100290 : data_o = 32'h3f3d853a ;
			32'h00100294 : data_o = 32'h9793872a ;
			32'h00100298 : data_o = 32'h17c10024 ;
			32'h0010029c : data_o = 32'ha82397a2 ;
			32'h001002a0 : data_o = 32'h2783fce7 ;
			32'h001002a4 : data_o = 32'h0785fec4 ;
			32'h001002a8 : data_o = 32'hfef42623 ;
			32'h001002ac : data_o = 32'hfec42703 ;
			32'h001002b0 : data_o = 32'hfae3478d ;
			32'h001002b4 : data_o = 32'h4529f8e7 ;
			32'h001002b8 : data_o = 32'h222328e9 ;
			32'h001002bc : data_o = 32'ha86dfe04 ;
			32'h001002c0 : data_o = 32'hfe042423 ;
			32'h001002c4 : data_o = 32'h0513a871 ;
			32'h001002c8 : data_o = 32'h20e107c0 ;
			32'h001002cc : data_o = 32'hfe042023 ;
			32'h001002d0 : data_o = 32'h2703a89d ;
			32'h001002d4 : data_o = 32'h478dfe44 ;
			32'h001002d8 : data_o = 32'h02e7c863 ;
			32'h001002dc : data_o = 32'hfe842783 ;
			32'h001002e0 : data_o = 32'h078a0786 ;
			32'h001002e4 : data_o = 32'h97a217c1 ;
			32'h001002e8 : data_o = 32'hfd07a683 ;
			32'h001002ec : data_o = 32'hfe442783 ;
			32'h001002f0 : data_o = 32'h00379713 ;
			32'h001002f4 : data_o = 32'hfe042783 ;
			32'h001002f8 : data_o = 32'h85be97ba ;
			32'h001002fc : data_o = 32'h3ddd8536 ;
			32'h00100300 : data_o = 32'h853e87aa ;
			32'h00100304 : data_o = 32'ha8052079 ;
			32'h00100308 : data_o = 32'hfe842783 ;
			32'h0010030c : data_o = 32'h07850786 ;
			32'h00100310 : data_o = 32'h17c1078a ;
			32'h00100314 : data_o = 32'ha68397a2 ;
			32'h00100318 : data_o = 32'h2783fd07 ;
			32'h0010031c : data_o = 32'h17f1fe44 ;
			32'h00100320 : data_o = 32'h00379713 ;
			32'h00100324 : data_o = 32'hfe042783 ;
			32'h00100328 : data_o = 32'h85be97ba ;
			32'h0010032c : data_o = 32'h35d98536 ;
			32'h00100330 : data_o = 32'h853e87aa ;
			32'h00100334 : data_o = 32'h051328b9 ;
			32'h00100338 : data_o = 32'h28a107c0 ;
			32'h0010033c : data_o = 32'hfe042783 ;
			32'h00100340 : data_o = 32'h20230785 ;
			32'h00100344 : data_o = 32'h2703fef4 ;
			32'h00100348 : data_o = 32'h479dfe04 ;
			32'h0010034c : data_o = 32'hf8e7d3e3 ;
			32'h00100350 : data_o = 32'h02000513 ;
			32'h00100354 : data_o = 32'h2783283d ;
			32'h00100358 : data_o = 32'h0785fe84 ;
			32'h0010035c : data_o = 32'hfef42423 ;
			32'h00100360 : data_o = 32'hfe842703 ;
			32'h00100364 : data_o = 32'hd0e3478d ;
			32'h00100368 : data_o = 32'h4529f6e7 ;
			32'h0010036c : data_o = 32'h2783201d ;
			32'h00100370 : data_o = 32'h0785fe44 ;
			32'h00100374 : data_o = 32'hfef42223 ;
			32'h00100378 : data_o = 32'hfe442703 ;
			32'h0010037c : data_o = 32'hd1e3479d ;
			32'h00100380 : data_o = 32'h4529f4e7 ;
			32'h00100384 : data_o = 32'h00012039 ;
			32'h00100388 : data_o = 32'h442640b6 ;
			32'h0010038c : data_o = 32'h61614496 ;
			32'h00100390 : data_o = 32'h11018082 ;
			32'h00100394 : data_o = 32'hcc22ce06 ;
			32'h00100398 : data_o = 32'h87aa1000 ;
			32'h0010039c : data_o = 32'hfef407a3 ;
			32'h001003a0 : data_o = 32'hfef44703 ;
			32'h001003a4 : data_o = 32'h166347a9 ;
			32'h001003a8 : data_o = 32'h45b500f7 ;
			32'h001003ac : data_o = 32'h80001537 ;
			32'h001003b0 : data_o = 32'h47832e2d ;
			32'h001003b4 : data_o = 32'h85befef4 ;
			32'h001003b8 : data_o = 32'h80001537 ;
			32'h001003bc : data_o = 32'h4783263d ;
			32'h001003c0 : data_o = 32'h853efef4 ;
			32'h001003c4 : data_o = 32'h446240f2 ;
			32'h001003c8 : data_o = 32'h80826105 ;
			32'h001003cc : data_o = 32'hc6061141 ;
			32'h001003d0 : data_o = 32'h0800c422 ;
			32'h001003d4 : data_o = 32'h80001537 ;
			32'h001003d8 : data_o = 32'h87aa24c5 ;
			32'h001003dc : data_o = 32'h40b2853e ;
			32'h001003e0 : data_o = 32'h01414422 ;
			32'h001003e4 : data_o = 32'h11018082 ;
			32'h001003e8 : data_o = 32'hcc22ce06 ;
			32'h001003ec : data_o = 32'h26231000 ;
			32'h001003f0 : data_o = 32'ha819fea4 ;
			32'h001003f4 : data_o = 32'hfec42783 ;
			32'h001003f8 : data_o = 32'h00178713 ;
			32'h001003fc : data_o = 32'hfee42623 ;
			32'h00100400 : data_o = 32'h0007c783 ;
			32'h00100404 : data_o = 32'h3771853e ;
			32'h00100408 : data_o = 32'hfec42783 ;
			32'h0010040c : data_o = 32'h0007c783 ;
			32'h00100410 : data_o = 32'h4781f3f5 ;
			32'h00100414 : data_o = 32'h40f2853e ;
			32'h00100418 : data_o = 32'h61054462 ;
			32'h0010041c : data_o = 32'h71798082 ;
			32'h00100420 : data_o = 32'hd422d606 ;
			32'h00100424 : data_o = 32'h2e231800 ;
			32'h00100428 : data_o = 32'h2623fca4 ;
			32'h0010042c : data_o = 32'ha891fe04 ;
			32'h00100430 : data_o = 32'hfdc42783 ;
			32'h00100434 : data_o = 32'h242383f1 ;
			32'h00100438 : data_o = 32'h2703fef4 ;
			32'h0010043c : data_o = 32'h47a5fe84 ;
			32'h00100440 : data_o = 32'h00e7cd63 ;
			32'h00100444 : data_o = 32'hfe842783 ;
			32'h00100448 : data_o = 32'h0ff7f793 ;
			32'h0010044c : data_o = 32'h03078793 ;
			32'h00100450 : data_o = 32'h0ff7f793 ;
			32'h00100454 : data_o = 32'h3f35853e ;
			32'h00100458 : data_o = 32'h2783a819 ;
			32'h0010045c : data_o = 32'hf793fe84 ;
			32'h00100460 : data_o = 32'h87930ff7 ;
			32'h00100464 : data_o = 32'hf7930377 ;
			32'h00100468 : data_o = 32'h853e0ff7 ;
			32'h0010046c : data_o = 32'h2783371d ;
			32'h00100470 : data_o = 32'h0792fdc4 ;
			32'h00100474 : data_o = 32'hfcf42e23 ;
			32'h00100478 : data_o = 32'hfec42783 ;
			32'h0010047c : data_o = 32'h26230785 ;
			32'h00100480 : data_o = 32'h2703fef4 ;
			32'h00100484 : data_o = 32'h479dfec4 ;
			32'h00100488 : data_o = 32'hfae7d4e3 ;
			32'h0010048c : data_o = 32'h00010001 ;
			32'h00100490 : data_o = 32'h542250b2 ;
			32'h00100494 : data_o = 32'h80826145 ;
			32'h00100498 : data_o = 32'hc6221141 ;
			32'h0010049c : data_o = 32'h07b70800 ;
			32'h001004a0 : data_o = 32'h07a10002 ;
			32'h001004a4 : data_o = 32'hc3984705 ;
			32'h001004a8 : data_o = 32'h44320001 ;
			32'h001004ac : data_o = 32'h80820141 ;
			32'h001004b0 : data_o = 32'hce221101 ;
			32'h001004b4 : data_o = 32'h27f31000 ;
			32'h001004b8 : data_o = 32'h26233410 ;
			32'h001004bc : data_o = 32'h2783fef4 ;
			32'h001004c0 : data_o = 32'h853efec4 ;
			32'h001004c4 : data_o = 32'h61054472 ;
			32'h001004c8 : data_o = 32'h11018082 ;
			32'h001004cc : data_o = 32'h1000ce22 ;
			32'h001004d0 : data_o = 32'h342027f3 ;
			32'h001004d4 : data_o = 32'hfef42623 ;
			32'h001004d8 : data_o = 32'hfec42783 ;
			32'h001004dc : data_o = 32'h4472853e ;
			32'h001004e0 : data_o = 32'h80826105 ;
			32'h001004e4 : data_o = 32'hce221101 ;
			32'h001004e8 : data_o = 32'h27f31000 ;
			32'h001004ec : data_o = 32'h26233430 ;
			32'h001004f0 : data_o = 32'h2783fef4 ;
			32'h001004f4 : data_o = 32'h853efec4 ;
			32'h001004f8 : data_o = 32'h61054472 ;
			32'h001004fc : data_o = 32'h11018082 ;
			32'h00100500 : data_o = 32'h1000ce22 ;
			32'h00100504 : data_o = 32'hb00027f3 ;
			32'h00100508 : data_o = 32'hfef42623 ;
			32'h0010050c : data_o = 32'hfec42783 ;
			32'h00100510 : data_o = 32'h4472853e ;
			32'h00100514 : data_o = 32'h80826105 ;
			32'h00100518 : data_o = 32'hc6221141 ;
			32'h0010051c : data_o = 32'h10730800 ;
			32'h00100520 : data_o = 32'h0001b000 ;
			32'h00100524 : data_o = 32'h01414432 ;
			32'h00100528 : data_o = 32'h71798082 ;
			32'h0010052c : data_o = 32'h1800d622 ;
			32'h00100530 : data_o = 32'hfca42e23 ;
			32'h00100534 : data_o = 32'hfcb42c23 ;
			32'h00100538 : data_o = 32'hfdc42703 ;
			32'h0010053c : data_o = 32'hf46347fd ;
			32'h00100540 : data_o = 32'h478500e7 ;
			32'h00100544 : data_o = 32'h0797a879 ;
			32'h00100548 : data_o = 32'h87930010 ;
			32'h0010054c : data_o = 32'h4398aba7 ;
			32'h00100550 : data_o = 32'hfdc42783 ;
			32'h00100554 : data_o = 32'h97ba078a ;
			32'h00100558 : data_o = 32'hfef42623 ;
			32'h0010055c : data_o = 32'hfd842703 ;
			32'h00100560 : data_o = 32'hfec42783 ;
			32'h00100564 : data_o = 32'h40f707b3 ;
			32'h00100568 : data_o = 32'hfef42423 ;
			32'h0010056c : data_o = 32'hfe842703 ;
			32'h00100570 : data_o = 32'h000807b7 ;
			32'h00100574 : data_o = 32'h00f75863 ;
			32'h00100578 : data_o = 32'hfe842703 ;
			32'h0010057c : data_o = 32'hfff807b7 ;
			32'h00100580 : data_o = 32'h00f75463 ;
			32'h00100584 : data_o = 32'ha8b14789 ;
			32'h00100588 : data_o = 32'hfe842783 ;
			32'h0010058c : data_o = 32'hfef42223 ;
			32'h00100590 : data_o = 32'hfe442783 ;
			32'h00100594 : data_o = 32'h01479713 ;
			32'h00100598 : data_o = 32'h7fe007b7 ;
			32'h0010059c : data_o = 32'h27838f7d ;
			32'h001005a0 : data_o = 32'h9693fe44 ;
			32'h001005a4 : data_o = 32'h07b70097 ;
			32'h001005a8 : data_o = 32'h8ff50010 ;
			32'h001005ac : data_o = 32'h26838f5d ;
			32'h001005b0 : data_o = 32'hf7b7fe44 ;
			32'h001005b4 : data_o = 32'h8ff5000f ;
			32'h001005b8 : data_o = 32'h27838f5d ;
			32'h001005bc : data_o = 32'h9693fe44 ;
			32'h001005c0 : data_o = 32'h07b700b7 ;
			32'h001005c4 : data_o = 32'h8ff58000 ;
			32'h001005c8 : data_o = 32'he7938fd9 ;
			32'h001005cc : data_o = 32'h202306f7 ;
			32'h001005d0 : data_o = 32'h2783fef4 ;
			32'h001005d4 : data_o = 32'h2703fec4 ;
			32'h001005d8 : data_o = 32'hc398fe04 ;
			32'h001005dc : data_o = 32'h0000100f ;
			32'h001005e0 : data_o = 32'h853e4781 ;
			32'h001005e4 : data_o = 32'h61455432 ;
			32'h001005e8 : data_o = 32'h11018082 ;
			32'h001005ec : data_o = 32'h1000ce22 ;
			32'h001005f0 : data_o = 32'hfea42623 ;
			32'h001005f4 : data_o = 32'hfec42783 ;
			32'h001005f8 : data_o = 32'h3047a073 ;
			32'h001005fc : data_o = 32'h44720001 ;
			32'h00100600 : data_o = 32'h80826105 ;
			32'h00100604 : data_o = 32'hce221101 ;
			32'h00100608 : data_o = 32'h26231000 ;
			32'h0010060c : data_o = 32'h2783fea4 ;
			32'h00100610 : data_o = 32'hb073fec4 ;
			32'h00100614 : data_o = 32'h00013047 ;
			32'h00100618 : data_o = 32'h61054472 ;
			32'h0010061c : data_o = 32'h11018082 ;
			32'h00100620 : data_o = 32'h1000ce22 ;
			32'h00100624 : data_o = 32'hfea42623 ;
			32'h00100628 : data_o = 32'hfec42783 ;
			32'h0010062c : data_o = 32'h47a1c789 ;
			32'h00100630 : data_o = 32'h3007a073 ;
			32'h00100634 : data_o = 32'h47a1a021 ;
			32'h00100638 : data_o = 32'h3007b073 ;
			32'h0010063c : data_o = 32'h44720001 ;
			32'h00100640 : data_o = 32'h80826105 ;
			32'h00100644 : data_o = 32'hc6061141 ;
			32'h00100648 : data_o = 32'h0800c422 ;
			32'h0010064c : data_o = 32'h00000517 ;
			32'h00100650 : data_o = 32'h68450513 ;
			32'h00100654 : data_o = 32'h05173b49 ;
			32'h00100658 : data_o = 32'h05130000 ;
			32'h0010065c : data_o = 32'h336168a5 ;
			32'h00100660 : data_o = 32'h00000517 ;
			32'h00100664 : data_o = 32'h69050513 ;
			32'h00100668 : data_o = 32'h35993bbd ;
			32'h0010066c : data_o = 32'h853e87aa ;
			32'h00100670 : data_o = 32'h0517337d ;
			32'h00100674 : data_o = 32'h05130000 ;
			32'h00100678 : data_o = 32'h33b568a5 ;
			32'h0010067c : data_o = 32'h87aa35b9 ;
			32'h00100680 : data_o = 32'h3b71853e ;
			32'h00100684 : data_o = 32'h00000517 ;
			32'h00100688 : data_o = 32'h68450513 ;
			32'h0010068c : data_o = 32'h3d993ba9 ;
			32'h00100690 : data_o = 32'h853e87aa ;
			32'h00100694 : data_o = 32'h45293369 ;
			32'h00100698 : data_o = 32'h000139ed ;
			32'h0010069c : data_o = 32'h1141bffd ;
			32'h001006a0 : data_o = 32'hc422c606 ;
			32'h001006a4 : data_o = 32'h65410800 ;
			32'h001006a8 : data_o = 32'h45053789 ;
			32'h001006ac : data_o = 32'h00013f8d ;
			32'h001006b0 : data_o = 32'h442240b2 ;
			32'h001006b4 : data_o = 32'h80820141 ;
			32'h001006b8 : data_o = 32'hd6227179 ;
			32'h001006bc : data_o = 32'h2e231800 ;
			32'h001006c0 : data_o = 32'h57fdfca4 ;
			32'h001006c4 : data_o = 32'hfef42623 ;
			32'h001006c8 : data_o = 32'hfdc42783 ;
			32'h001006cc : data_o = 32'h439c07a1 ;
			32'h001006d0 : data_o = 32'he7918b85 ;
			32'h001006d4 : data_o = 32'hfdc42783 ;
			32'h001006d8 : data_o = 32'h2623439c ;
			32'h001006dc : data_o = 32'h2783fef4 ;
			32'h001006e0 : data_o = 32'h853efec4 ;
			32'h001006e4 : data_o = 32'h61455432 ;
			32'h001006e8 : data_o = 32'h11018082 ;
			32'h001006ec : data_o = 32'h1000ce22 ;
			32'h001006f0 : data_o = 32'hfea42623 ;
			32'h001006f4 : data_o = 32'h05a387ae ;
			32'h001006f8 : data_o = 32'h0001fef4 ;
			32'h001006fc : data_o = 32'hfec42783 ;
			32'h00100700 : data_o = 32'h439c07a1 ;
			32'h00100704 : data_o = 32'hfbfd8b89 ;
			32'h00100708 : data_o = 32'hfec42783 ;
			32'h0010070c : data_o = 32'h47030791 ;
			32'h00100710 : data_o = 32'hc398feb4 ;
			32'h00100714 : data_o = 32'h44720001 ;
			32'h00100718 : data_o = 32'h80826105 ;
			32'h0010071c : data_o = 32'hce221101 ;
			32'h00100720 : data_o = 32'h24231000 ;
			32'h00100724 : data_o = 32'h2623fea4 ;
			32'h00100728 : data_o = 32'h26b7feb4 ;
			32'h0010072c : data_o = 32'h06a10800 ;
			32'h00100730 : data_o = 32'hc290567d ;
			32'h00100734 : data_o = 32'hfec42683 ;
			32'h00100738 : data_o = 32'h0006d713 ;
			32'h0010073c : data_o = 32'h26b74781 ;
			32'h00100740 : data_o = 32'h06b10800 ;
			32'h00100744 : data_o = 32'hc29c87ba ;
			32'h00100748 : data_o = 32'h080027b7 ;
			32'h0010074c : data_o = 32'h270307a1 ;
			32'h00100750 : data_o = 32'hc398fe84 ;
			32'h00100754 : data_o = 32'h44720001 ;
			32'h00100758 : data_o = 32'h80826105 ;
			32'h0010075c : data_o = 32'hd6067179 ;
			32'h00100760 : data_o = 32'h1800d422 ;
			32'h00100764 : data_o = 32'hfca42c23 ;
			32'h00100768 : data_o = 32'hfcb42e23 ;
			32'h0010076c : data_o = 32'h242320fd ;
			32'h00100770 : data_o = 32'h2623fea4 ;
			32'h00100774 : data_o = 32'h2603feb4 ;
			32'h00100778 : data_o = 32'h2683fe84 ;
			32'h0010077c : data_o = 32'h2503fec4 ;
			32'h00100780 : data_o = 32'h2583fd84 ;
			32'h00100784 : data_o = 32'h0733fdc4 ;
			32'h00100788 : data_o = 32'h883a00a6 ;
			32'h0010078c : data_o = 32'h00c83833 ;
			32'h00100790 : data_o = 32'h00b687b3 ;
			32'h00100794 : data_o = 32'h00f806b3 ;
			32'h00100798 : data_o = 32'h242387b6 ;
			32'h0010079c : data_o = 32'h2623fee4 ;
			32'h001007a0 : data_o = 32'h2503fef4 ;
			32'h001007a4 : data_o = 32'h2583fe84 ;
			32'h001007a8 : data_o = 32'h3f8dfec4 ;
			32'h001007ac : data_o = 32'h50b20001 ;
			32'h001007b0 : data_o = 32'h61455422 ;
			32'h001007b4 : data_o = 32'h715d8082 ;
			32'h001007b8 : data_o = 32'hc496c686 ;
			32'h001007bc : data_o = 32'hc09ec29a ;
			32'h001007c0 : data_o = 32'hdc2ade22 ;
			32'h001007c4 : data_o = 32'hd832da2e ;
			32'h001007c8 : data_o = 32'hd43ad636 ;
			32'h001007cc : data_o = 32'hd042d23e ;
			32'h001007d0 : data_o = 32'hcc72ce46 ;
			32'h001007d4 : data_o = 32'hc87aca76 ;
			32'h001007d8 : data_o = 32'h0880c67e ;
			32'h001007dc : data_o = 32'h00100797 ;
			32'h001007e0 : data_o = 32'h83c78793 ;
			32'h001007e4 : data_o = 32'h43dc4398 ;
			32'h001007e8 : data_o = 32'h85be853a ;
			32'h001007ec : data_o = 32'h07973f85 ;
			32'h001007f0 : data_o = 32'h87930010 ;
			32'h001007f4 : data_o = 32'h43988227 ;
			32'h001007f8 : data_o = 32'h450543dc ;
			32'h001007fc : data_o = 32'h06334581 ;
			32'h00100800 : data_o = 32'h883200a7 ;
			32'h00100804 : data_o = 32'h00e83833 ;
			32'h00100808 : data_o = 32'h00b786b3 ;
			32'h0010080c : data_o = 32'h00d807b3 ;
			32'h00100810 : data_o = 32'h873286be ;
			32'h00100814 : data_o = 32'hf69787b6 ;
			32'h00100818 : data_o = 32'h8693000f ;
			32'h0010081c : data_o = 32'hc2987fa6 ;
			32'h00100820 : data_o = 32'h0001c2dc ;
			32'h00100824 : data_o = 32'h42a640b6 ;
			32'h00100828 : data_o = 32'h43864316 ;
			32'h0010082c : data_o = 32'h55625472 ;
			32'h00100830 : data_o = 32'h564255d2 ;
			32'h00100834 : data_o = 32'h572256b2 ;
			32'h00100838 : data_o = 32'h58025792 ;
			32'h0010083c : data_o = 32'h4e6248f2 ;
			32'h00100840 : data_o = 32'h4f424ed2 ;
			32'h00100844 : data_o = 32'h61614fb2 ;
			32'h00100848 : data_o = 32'h30200073 ;
			32'h0010084c : data_o = 32'hc6221141 ;
			32'h00100850 : data_o = 32'h00010800 ;
			32'h00100854 : data_o = 32'h01414432 ;
			32'h00100858 : data_o = 32'h11018082 ;
			32'h0010085c : data_o = 32'h1000ce22 ;
			32'h00100860 : data_o = 32'h08002837 ;
			32'h00100864 : data_o = 32'h28030811 ;
			32'h00100868 : data_o = 32'h26230008 ;
			32'h0010086c : data_o = 32'h2837ff04 ;
			32'h00100870 : data_o = 32'h28030800 ;
			32'h00100874 : data_o = 32'h24230008 ;
			32'h00100878 : data_o = 32'h2837ff04 ;
			32'h0010087c : data_o = 32'h08110800 ;
			32'h00100880 : data_o = 32'h00082803 ;
			32'h00100884 : data_o = 32'hfec42883 ;
			32'h00100888 : data_o = 32'hfd089ce3 ;
			32'h0010088c : data_o = 32'hfec42803 ;
			32'h00100890 : data_o = 32'h45818542 ;
			32'h00100894 : data_o = 32'h00051793 ;
			32'h00100898 : data_o = 32'h25834701 ;
			32'h0010089c : data_o = 32'h862efe84 ;
			32'h001008a0 : data_o = 32'h65b34681 ;
			32'h001008a4 : data_o = 32'h202300c7 ;
			32'h001008a8 : data_o = 32'h8fd5feb4 ;
			32'h001008ac : data_o = 32'hfef42223 ;
			32'h001008b0 : data_o = 32'hfe042703 ;
			32'h001008b4 : data_o = 32'hfe442783 ;
			32'h001008b8 : data_o = 32'h85be853a ;
			32'h001008bc : data_o = 32'h61054472 ;
			32'h001008c0 : data_o = 32'h11418082 ;
			32'h001008c4 : data_o = 32'h0800c622 ;
			32'h001008c8 : data_o = 32'h000ff797 ;
			32'h001008cc : data_o = 32'h74878793 ;
			32'h001008d0 : data_o = 32'h43dc4398 ;
			32'h001008d4 : data_o = 32'h85be853a ;
			32'h001008d8 : data_o = 32'h01414432 ;
			32'h001008dc : data_o = 32'h11018082 ;
			32'h001008e0 : data_o = 32'hcc22ce06 ;
			32'h001008e4 : data_o = 32'h24231000 ;
			32'h001008e8 : data_o = 32'h2623fea4 ;
			32'h001008ec : data_o = 32'hf797feb4 ;
			32'h001008f0 : data_o = 32'h8793000f ;
			32'h001008f4 : data_o = 32'h46817227 ;
			32'h001008f8 : data_o = 32'hc3944701 ;
			32'h001008fc : data_o = 32'hf697c3d8 ;
			32'h00100900 : data_o = 32'h8693000f ;
			32'h00100904 : data_o = 32'h270371a6 ;
			32'h00100908 : data_o = 32'h2783fe84 ;
			32'h0010090c : data_o = 32'hc298fec4 ;
			32'h00100910 : data_o = 32'h2503c2dc ;
			32'h00100914 : data_o = 32'h2583fe84 ;
			32'h00100918 : data_o = 32'h3589fec4 ;
			32'h0010091c : data_o = 32'h08000513 ;
			32'h00100920 : data_o = 32'h450531e9 ;
			32'h00100924 : data_o = 32'h000139ed ;
			32'h00100928 : data_o = 32'h446240f2 ;
			32'h0010092c : data_o = 32'h80826105 ;
			32'h00100930 : data_o = 32'hc6221141 ;
			32'h00100934 : data_o = 32'h07930800 ;
			32'h00100938 : data_o = 32'hb0730800 ;
			32'h0010093c : data_o = 32'h00013047 ;
			32'h00100940 : data_o = 32'h01414432 ;
			32'h00100944 : data_o = 32'h11018082 ;
			32'h00100948 : data_o = 32'h1000ce22 ;
			32'h0010094c : data_o = 32'hfea42623 ;
			32'h00100950 : data_o = 32'hfeb42423 ;
			32'h00100954 : data_o = 32'hfec42783 ;
			32'h00100958 : data_o = 32'hfe842703 ;
			32'h0010095c : data_o = 32'h0001c398 ;
			32'h00100960 : data_o = 32'h61054472 ;
			32'h00100964 : data_o = 32'h11018082 ;
			32'h00100968 : data_o = 32'h1000ce22 ;
			32'h0010096c : data_o = 32'hfea42623 ;
			32'h00100970 : data_o = 32'hfec42783 ;
			32'h00100974 : data_o = 32'h853e439c ;
			32'h00100978 : data_o = 32'h61054472 ;
			32'h0010097c : data_o = 32'h71798082 ;
			32'h00100980 : data_o = 32'hd422d606 ;
			32'h00100984 : data_o = 32'h2e231800 ;
			32'h00100988 : data_o = 32'h2c23fca4 ;
			32'h0010098c : data_o = 32'h2a23fcb4 ;
			32'h00100990 : data_o = 32'h2503fcc4 ;
			32'h00100994 : data_o = 32'h3fc1fdc4 ;
			32'h00100998 : data_o = 32'hfea42623 ;
			32'h0010099c : data_o = 32'hfd842783 ;
			32'h001009a0 : data_o = 32'h17b34705 ;
			32'h001009a4 : data_o = 32'hc79300f7 ;
			32'h001009a8 : data_o = 32'h873efff7 ;
			32'h001009ac : data_o = 32'hfec42783 ;
			32'h001009b0 : data_o = 32'h26238ff9 ;
			32'h001009b4 : data_o = 32'h2783fef4 ;
			32'h001009b8 : data_o = 32'h2703fd84 ;
			32'h001009bc : data_o = 32'h17b3fd44 ;
			32'h001009c0 : data_o = 32'h270300f7 ;
			32'h001009c4 : data_o = 32'h8fd9fec4 ;
			32'h001009c8 : data_o = 32'hfef42623 ;
			32'h001009cc : data_o = 32'hfec42583 ;
			32'h001009d0 : data_o = 32'hfdc42503 ;
			32'h001009d4 : data_o = 32'h00013f8d ;
			32'h001009d8 : data_o = 32'h542250b2 ;
			32'h001009dc : data_o = 32'h80826145 ;
			32'h001009e0 : data_o = 32'hd6067179 ;
			32'h001009e4 : data_o = 32'h1800d422 ;
			32'h001009e8 : data_o = 32'hfca42e23 ;
			32'h001009ec : data_o = 32'hfcb42c23 ;
			32'h001009f0 : data_o = 32'hfdc42503 ;
			32'h001009f4 : data_o = 32'h26233f8d ;
			32'h001009f8 : data_o = 32'h2783fea4 ;
			32'h001009fc : data_o = 32'h2703fd84 ;
			32'h00100a00 : data_o = 32'h57b3fec4 ;
			32'h00100a04 : data_o = 32'h8b8500f7 ;
			32'h00100a08 : data_o = 32'h50b2853e ;
			32'h00100a0c : data_o = 32'h61455422 ;
			32'h00100a10 : data_o = 32'h11018082 ;
			32'h00100a14 : data_o = 32'h1000ce22 ;
			32'h00100a18 : data_o = 32'hfea42623 ;
			32'h00100a1c : data_o = 32'h700007b7 ;
			32'h00100a20 : data_o = 32'h270307c1 ;
			32'h00100a24 : data_o = 32'hc398fec4 ;
			32'h00100a28 : data_o = 32'h44720001 ;
			32'h00100a2c : data_o = 32'h80826105 ;
			32'h00100a30 : data_o = 32'hd6227179 ;
			32'h00100a34 : data_o = 32'h2e231800 ;
			32'h00100a38 : data_o = 32'h2783fca4 ;
			32'h00100a3c : data_o = 32'hc783fdc4 ;
			32'h00100a40 : data_o = 32'h873e0007 ;
			32'h00100a44 : data_o = 32'hfdc42783 ;
			32'h00100a48 : data_o = 32'hc7830785 ;
			32'h00100a4c : data_o = 32'h07a20007 ;
			32'h00100a50 : data_o = 32'h27838f5d ;
			32'h00100a54 : data_o = 32'h0789fdc4 ;
			32'h00100a58 : data_o = 32'h0007c783 ;
			32'h00100a5c : data_o = 32'h8f5d07c2 ;
			32'h00100a60 : data_o = 32'hfdc42783 ;
			32'h00100a64 : data_o = 32'hc783078d ;
			32'h00100a68 : data_o = 32'h07e20007 ;
			32'h00100a6c : data_o = 32'h26238fd9 ;
			32'h00100a70 : data_o = 32'h07b7fef4 ;
			32'h00100a74 : data_o = 32'h07e17000 ;
			32'h00100a78 : data_o = 32'hfec42703 ;
			32'h00100a7c : data_o = 32'h0001c398 ;
			32'h00100a80 : data_o = 32'h61455432 ;
			32'h00100a84 : data_o = 32'h11418082 ;
			32'h00100a88 : data_o = 32'h0800c622 ;
			32'h00100a8c : data_o = 32'h700007b7 ;
			32'h00100a90 : data_o = 32'h02078793 ;
			32'h00100a94 : data_o = 32'hc3984705 ;
			32'h00100a98 : data_o = 32'h44320001 ;
			32'h00100a9c : data_o = 32'h80820141 ;
			32'h00100aa0 : data_o = 32'hc6221141 ;
			32'h00100aa4 : data_o = 32'h00010800 ;
			32'h00100aa8 : data_o = 32'h700007b7 ;
			32'h00100aac : data_o = 32'h02478793 ;
			32'h00100ab0 : data_o = 32'hdbfd439c ;
			32'h00100ab4 : data_o = 32'h700007b7 ;
			32'h00100ab8 : data_o = 32'h02878793 ;
			32'h00100abc : data_o = 32'h853e439c ;
			32'h00100ac0 : data_o = 32'h01414432 ;
			32'h00100ac4 : data_o = 32'h11418082 ;
			32'h00100ac8 : data_o = 32'hc422c606 ;
			32'h00100acc : data_o = 32'h05370800 ;
			32'h00100ad0 : data_o = 32'h3e210002 ;
			32'h00100ad4 : data_o = 32'h36a14505 ;
			32'h00100ad8 : data_o = 32'h700007b7 ;
			32'h00100adc : data_o = 32'h03078793 ;
			32'h00100ae0 : data_o = 32'hc3984705 ;
			32'h00100ae4 : data_o = 32'h40b20001 ;
			32'h00100ae8 : data_o = 32'h01414422 ;
			32'h00100aec : data_o = 32'h11418082 ;
			32'h00100af0 : data_o = 32'hc422c606 ;
			32'h00100af4 : data_o = 32'h07b70800 ;
			32'h00100af8 : data_o = 32'h87937000 ;
			32'h00100afc : data_o = 32'ha0230307 ;
			32'h00100b00 : data_o = 32'h05370007 ;
			32'h00100b04 : data_o = 32'h3cfd0002 ;
			32'h00100b08 : data_o = 32'h40b20001 ;
			32'h00100b0c : data_o = 32'h01414422 ;
			32'h00100b10 : data_o = 32'h11018082 ;
			32'h00100b14 : data_o = 32'h1000ce22 ;
			32'h00100b18 : data_o = 32'hfea42623 ;
			32'h00100b1c : data_o = 32'h700007b7 ;
			32'h00100b20 : data_o = 32'h03478793 ;
			32'h00100b24 : data_o = 32'hfec42703 ;
			32'h00100b28 : data_o = 32'h0001c398 ;
			32'h00100b2c : data_o = 32'h61054472 ;
			32'h00100b30 : data_o = 32'h11018082 ;
			32'h00100b34 : data_o = 32'h1000ce22 ;
			32'h00100b38 : data_o = 32'hfea42623 ;
			32'h00100b3c : data_o = 32'h700007b7 ;
			32'h00100b40 : data_o = 32'h03c78793 ;
			32'h00100b44 : data_o = 32'hfec40713 ;
			32'h00100b48 : data_o = 32'h0001c398 ;
			32'h00100b4c : data_o = 32'h61054472 ;
			32'h00100b50 : data_o = 32'h11018082 ;
			32'h00100b54 : data_o = 32'h1000ce22 ;
			32'h00100b58 : data_o = 32'hfea42623 ;
			32'h00100b5c : data_o = 32'h700007b7 ;
			32'h00100b60 : data_o = 32'h03878793 ;
			32'h00100b64 : data_o = 32'hfec42703 ;
			32'h00100b68 : data_o = 32'h0001c398 ;
			32'h00100b6c : data_o = 32'h61054472 ;
			32'h00100b70 : data_o = 32'h11418082 ;
			32'h00100b74 : data_o = 32'h0800c622 ;
			32'h00100b78 : data_o = 32'h700007b7 ;
			32'h00100b7c : data_o = 32'h04078793 ;
			32'h00100b80 : data_o = 32'hf793439c ;
			32'h00100b84 : data_o = 32'h853e0ff7 ;
			32'h00100b88 : data_o = 32'h01414432 ;
			32'h00100b8c : data_o = 32'h11418082 ;
			32'h00100b90 : data_o = 32'h0800c622 ;
			32'h00100b94 : data_o = 32'h700007b7 ;
			32'h00100b98 : data_o = 32'h04478793 ;
			32'h00100b9c : data_o = 32'hc3984705 ;
			32'h00100ba0 : data_o = 32'h44320001 ;
			32'h00100ba4 : data_o = 32'h80820141 ;
			32'h00100ba8 : data_o = 32'hc6221141 ;
			32'h00100bac : data_o = 32'h07b70800 ;
			32'h00100bb0 : data_o = 32'h87937000 ;
			32'h00100bb4 : data_o = 32'ha0230447 ;
			32'h00100bb8 : data_o = 32'h00010007 ;
			32'h00100bbc : data_o = 32'h01414432 ;
			32'h00100bc0 : data_o = 32'h11018082 ;
			32'h00100bc4 : data_o = 32'h1000ce22 ;
			32'h00100bc8 : data_o = 32'hfea42623 ;
			32'h00100bcc : data_o = 32'h700007b7 ;
			32'h00100bd0 : data_o = 32'h04878793 ;
			32'h00100bd4 : data_o = 32'hfec42703 ;
			32'h00100bd8 : data_o = 32'h0001c398 ;
			32'h00100bdc : data_o = 32'h61054472 ;
			32'h00100be0 : data_o = 32'h11018082 ;
			32'h00100be4 : data_o = 32'h1000ce22 ;
			32'h00100be8 : data_o = 32'hfea42623 ;
			32'h00100bec : data_o = 32'h700007b7 ;
			32'h00100bf0 : data_o = 32'h04c78793 ;
			32'h00100bf4 : data_o = 32'hfec42703 ;
			32'h00100bf8 : data_o = 32'h0001c398 ;
			32'h00100bfc : data_o = 32'h61054472 ;
			32'h00100c00 : data_o = 32'h11018082 ;
			32'h00100c04 : data_o = 32'h1000ce22 ;
			32'h00100c08 : data_o = 32'hfea42623 ;
			32'h00100c0c : data_o = 32'h873287ae ;
			32'h00100c10 : data_o = 32'hfef405a3 ;
			32'h00100c14 : data_o = 32'h052387ba ;
			32'h00100c18 : data_o = 32'h2783fef4 ;
			32'h00100c1c : data_o = 32'h439cfec4 ;
			32'h00100c20 : data_o = 32'hfeb44703 ;
			32'h00100c24 : data_o = 32'h7693070e ;
			32'h00100c28 : data_o = 32'h17370187 ;
			32'h00100c2c : data_o = 32'h07137000 ;
			32'h00100c30 : data_o = 32'h8ed98007 ;
			32'h00100c34 : data_o = 32'hfea44703 ;
			32'h00100c38 : data_o = 32'h8f558b15 ;
			32'h00100c3c : data_o = 32'hfff7c793 ;
			32'h00100c40 : data_o = 32'h0001c31c ;
			32'h00100c44 : data_o = 32'h61054472 ;
			32'h00100c48 : data_o = 32'hf06f8082 ;
			32'h00100c4c : data_o = 32'h00939fbf ;
			32'h00100c50 : data_o = 32'h81060000 ;
			32'h00100c54 : data_o = 32'h82068186 ;
			32'h00100c58 : data_o = 32'h83068286 ;
			32'h00100c5c : data_o = 32'h84068386 ;
			32'h00100c60 : data_o = 32'h85068486 ;
			32'h00100c64 : data_o = 32'h86068586 ;
			32'h00100c68 : data_o = 32'h87068686 ;
			32'h00100c6c : data_o = 32'h88068786 ;
			32'h00100c70 : data_o = 32'h89068886 ;
			32'h00100c74 : data_o = 32'h8a068986 ;
			32'h00100c78 : data_o = 32'h8b068a86 ;
			32'h00100c7c : data_o = 32'h8c068b86 ;
			32'h00100c80 : data_o = 32'h8d068c86 ;
			32'h00100c84 : data_o = 32'h8e068d86 ;
			32'h00100c88 : data_o = 32'h8f068e86 ;
			32'h00100c8c : data_o = 32'hf1178f86 ;
			32'h00100c90 : data_o = 32'h01130010 ;
			32'h00100c94 : data_o = 32'hfd173721 ;
			32'h00100c98 : data_o = 32'h0d13000f ;
			32'h00100c9c : data_o = 32'hfd97372d ;
			32'h00100ca0 : data_o = 32'h8d93000f ;
			32'h00100ca4 : data_o = 32'h5763382d ;
			32'h00100ca8 : data_o = 32'h202301bd ;
			32'h00100cac : data_o = 32'h0d11000d ;
			32'h00100cb0 : data_o = 32'hffaddde3 ;
			32'h00100cb4 : data_o = 32'h45814501 ;
			32'h00100cb8 : data_o = 32'hc38ff0ef ;
			32'h00100cbc : data_o = 32'h000202b7 ;
			32'h00100cc0 : data_o = 32'h430502a1 ;
			32'h00100cc4 : data_o = 32'h0062a023 ;
			32'h00100cc8 : data_o = 32'h10500073 ;
			32'h00100ccc : data_o = 32'h0000bff5 ;
			32'h00100cd0 : data_o = 32'h45435845 ;
			32'h00100cd4 : data_o = 32'h4f495450 ;
			32'h00100cd8 : data_o = 32'h2121214e ;
			32'h00100cdc : data_o = 32'h0000000a ;
			32'h00100ce0 : data_o = 32'h3d3d3d3d ;
			32'h00100ce4 : data_o = 32'h3d3d3d3d ;
			32'h00100ce8 : data_o = 32'h3d3d3d3d ;
			32'h00100cec : data_o = 32'h0000000a ;
			32'h00100cf0 : data_o = 32'h4350454d ;
			32'h00100cf4 : data_o = 32'h2020203a ;
			32'h00100cf8 : data_o = 32'h00007830 ;
			32'h00100cfc : data_o = 32'h41434d0a ;
			32'h00100d00 : data_o = 32'h3a455355 ;
			32'h00100d04 : data_o = 32'h00783020 ;
			32'h00100d08 : data_o = 32'h56544d0a ;
			32'h00100d0c : data_o = 32'h203a4c41 ;
			32'h00100d10 : data_o = 32'h00783020 ;
			32'h00100d14 : data_o = 32'h00100000 ;
			default : data_o = 32'h00000000 ;
		endcase 
	end
endmodule
