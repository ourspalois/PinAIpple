module rom_1p #(
	int Depth, 
 	int DATA_WIDTH = 32, 
 	int ADDR_WIDTH = 32 
 ) (
	input logic clk_i, 
	input logic req_i, 
	input logic [ADDR_WIDTH-1:0] addr_i, 
	output logic [DATA_WIDTH-1:0] data_o 
 );
	always_ff @(posedge clk_i) begin
		case (addr_i)
			32'h00100000 : data_o = 32'h2c00006f ;
			32'h00100004 : data_o = 32'h2bc0006f ;
			32'h00100008 : data_o = 32'h2b80006f ;
			32'h0010000c : data_o = 32'h2b40006f ;
			32'h00100010 : data_o = 32'h2b00006f ;
			32'h00100014 : data_o = 32'h2ac0006f ;
			32'h00100018 : data_o = 32'h2a80006f ;
			32'h0010001c : data_o = 32'h2a40006f ;
			32'h00100020 : data_o = 32'h2a00006f ;
			32'h00100024 : data_o = 32'h29c0006f ;
			32'h00100028 : data_o = 32'h2980006f ;
			32'h0010002c : data_o = 32'h2940006f ;
			32'h00100030 : data_o = 32'h2900006f ;
			32'h00100034 : data_o = 32'h28c0006f ;
			32'h00100038 : data_o = 32'h2880006f ;
			32'h0010003c : data_o = 32'h2840006f ;
			32'h00100040 : data_o = 32'h2800006f ;
			32'h00100044 : data_o = 32'h06c0006f ;
			32'h00100048 : data_o = 32'h2780006f ;
			32'h0010004c : data_o = 32'h2740006f ;
			32'h00100050 : data_o = 32'h2700006f ;
			32'h00100054 : data_o = 32'h26c0006f ;
			32'h00100058 : data_o = 32'h2680006f ;
			32'h0010005c : data_o = 32'h2640006f ;
			32'h00100060 : data_o = 32'h2600006f ;
			32'h00100064 : data_o = 32'h25c0006f ;
			32'h00100068 : data_o = 32'h2580006f ;
			32'h0010006c : data_o = 32'h2540006f ;
			32'h00100070 : data_o = 32'h2500006f ;
			32'h00100074 : data_o = 32'h24c0006f ;
			32'h00100078 : data_o = 32'h2480006f ;
			32'h0010007c : data_o = 32'h2440006f ;
			32'h00100080 : data_o = 32'h4d20006f ;
			32'h00100084 : data_o = 32'h08134781 ;
			32'h00100088 : data_o = 32'h06130300 ;
			32'h0010008c : data_o = 32'h06930310 ;
			32'h00100090 : data_o = 32'ha0390200 ;
			32'h00100094 : data_o = 32'h01058023 ;
			32'h00100098 : data_o = 32'h05850785 ;
			32'h0010009c : data_o = 32'h00d78963 ;
			32'h001000a0 : data_o = 32'h00f55733 ;
			32'h001000a4 : data_o = 32'hd77d8b05 ;
			32'h001000a8 : data_o = 32'h00c58023 ;
			32'h001000ac : data_o = 32'h8082b7f5 ;
			32'h001000b0 : data_o = 32'hde067139 ;
			32'h001000b4 : data_o = 32'hda1adc16 ;
			32'h001000b8 : data_o = 32'hd62ad81e ;
			32'h001000bc : data_o = 32'hd232d42e ;
			32'h001000c0 : data_o = 32'hce3ad036 ;
			32'h001000c4 : data_o = 32'hca42cc3e ;
			32'h001000c8 : data_o = 32'hc672c846 ;
			32'h001000cc : data_o = 32'hc27ac476 ;
			32'h001000d0 : data_o = 32'h26f9c07e ;
			32'h001000d4 : data_o = 32'h00100797 ;
			32'h001000d8 : data_o = 32'hf2a7ac23 ;
			32'h001000dc : data_o = 32'h07174785 ;
			32'h001000e0 : data_o = 32'h25230010 ;
			32'h001000e4 : data_o = 32'h50f2f2f7 ;
			32'h001000e8 : data_o = 32'h535252e2 ;
			32'h001000ec : data_o = 32'h553253c2 ;
			32'h001000f0 : data_o = 32'h561255a2 ;
			32'h001000f4 : data_o = 32'h47725682 ;
			32'h001000f8 : data_o = 32'h485247e2 ;
			32'h001000fc : data_o = 32'h4e3248c2 ;
			32'h00100100 : data_o = 32'h4f124ea2 ;
			32'h00100104 : data_o = 32'h61214f82 ;
			32'h00100108 : data_o = 32'h30200073 ;
			32'h0010010c : data_o = 32'hc6061141 ;
			32'h00100110 : data_o = 32'h0413c422 ;
			32'h00100114 : data_o = 32'h28690fd0 ;
			32'h00100118 : data_o = 32'h0ff57513 ;
			32'h0010011c : data_o = 32'hfff50793 ;
			32'h00100120 : data_o = 32'h0ff7f793 ;
			32'h00100124 : data_o = 32'hfef469e3 ;
			32'h00100128 : data_o = 32'h442240b2 ;
			32'h0010012c : data_o = 32'h80820141 ;
			32'h00100130 : data_o = 32'hd6067179 ;
			32'h00100134 : data_o = 32'hd226d422 ;
			32'h00100138 : data_o = 32'h800007b7 ;
			32'h0010013c : data_o = 32'hc3984705 ;
			32'h00100140 : data_o = 32'h06100513 ;
			32'h00100144 : data_o = 32'h17b72089 ;
			32'h00100148 : data_o = 32'ha7037000 ;
			32'h0010014c : data_o = 32'h07978007 ;
			32'h00100150 : data_o = 32'h87930010 ;
			32'h00100154 : data_o = 32'hc398ebe7 ;
			32'h00100158 : data_o = 32'h858a4388 ;
			32'h0010015c : data_o = 32'h05133725 ;
			32'h00100160 : data_o = 32'h201507c0 ;
			32'h00100164 : data_o = 32'h1004840a ;
			32'h00100168 : data_o = 32'h00044503 ;
			32'h0010016c : data_o = 32'h05132829 ;
			32'h00100170 : data_o = 32'h281107c0 ;
			32'h00100174 : data_o = 32'h19e30405 ;
			32'h00100178 : data_o = 32'h4501fe94 ;
			32'h0010017c : data_o = 32'h542250b2 ;
			32'h00100180 : data_o = 32'h61455492 ;
			32'h00100184 : data_o = 32'h11418082 ;
			32'h00100188 : data_o = 32'hc422c606 ;
			32'h0010018c : data_o = 32'h47a9842a ;
			32'h00100190 : data_o = 32'h00f50b63 ;
			32'h00100194 : data_o = 32'h153785a2 ;
			32'h00100198 : data_o = 32'h2a518000 ;
			32'h0010019c : data_o = 32'h40b28522 ;
			32'h001001a0 : data_o = 32'h01414422 ;
			32'h001001a4 : data_o = 32'h45b58082 ;
			32'h001001a8 : data_o = 32'h80001537 ;
			32'h001001ac : data_o = 32'hb7dd2249 ;
			32'h001001b0 : data_o = 32'hc6061141 ;
			32'h001001b4 : data_o = 32'h80001537 ;
			32'h001001b8 : data_o = 32'h40b222a5 ;
			32'h001001bc : data_o = 32'h80820141 ;
			32'h001001c0 : data_o = 32'hc6061141 ;
			32'h001001c4 : data_o = 32'h842ac422 ;
			32'h001001c8 : data_o = 32'h00054503 ;
			32'h001001cc : data_o = 32'h0405c511 ;
			32'h001001d0 : data_o = 32'h45033f5d ;
			32'h001001d4 : data_o = 32'hfd650004 ;
			32'h001001d8 : data_o = 32'h40b24501 ;
			32'h001001dc : data_o = 32'h01414422 ;
			32'h001001e0 : data_o = 32'h11418082 ;
			32'h001001e4 : data_o = 32'hc422c606 ;
			32'h001001e8 : data_o = 32'hc04ac226 ;
			32'h001001ec : data_o = 32'h44a1842a ;
			32'h001001f0 : data_o = 32'ha0394925 ;
			32'h001001f4 : data_o = 32'h03750513 ;
			32'h001001f8 : data_o = 32'h04123779 ;
			32'h001001fc : data_o = 32'hc88914fd ;
			32'h00100200 : data_o = 32'h01c45513 ;
			32'h00100204 : data_o = 32'hfea948e3 ;
			32'h00100208 : data_o = 32'h03050513 ;
			32'h0010020c : data_o = 32'hb7f53fad ;
			32'h00100210 : data_o = 32'h442240b2 ;
			32'h00100214 : data_o = 32'h49024492 ;
			32'h00100218 : data_o = 32'h80820141 ;
			32'h0010021c : data_o = 32'h000207b7 ;
			32'h00100220 : data_o = 32'hc7984705 ;
			32'h00100224 : data_o = 32'h25738082 ;
			32'h00100228 : data_o = 32'h80823410 ;
			32'h0010022c : data_o = 32'h34202573 ;
			32'h00100230 : data_o = 32'h25738082 ;
			32'h00100234 : data_o = 32'h80823430 ;
			32'h00100238 : data_o = 32'hb0002573 ;
			32'h0010023c : data_o = 32'h10738082 ;
			32'h00100240 : data_o = 32'h8082b000 ;
			32'h00100244 : data_o = 32'hec6347fd ;
			32'h00100248 : data_o = 32'h050a04a7 ;
			32'h0010024c : data_o = 32'h00100717 ;
			32'h00100250 : data_o = 32'hdb472703 ;
			32'h00100254 : data_o = 32'h8d99972a ;
			32'h00100258 : data_o = 32'h000807b7 ;
			32'h0010025c : data_o = 32'h06b797ae ;
			32'h00100260 : data_o = 32'h45090010 ;
			32'h00100264 : data_o = 32'h02d7fe63 ;
			32'h00100268 : data_o = 32'h01459793 ;
			32'h0010026c : data_o = 32'h7fe006b7 ;
			32'h00100270 : data_o = 32'h96938ff5 ;
			32'h00100274 : data_o = 32'h063700b5 ;
			32'h00100278 : data_o = 32'h8ef18000 ;
			32'h0010027c : data_o = 32'hf6b78fd5 ;
			32'h00100280 : data_o = 32'h8eed000f ;
			32'h00100284 : data_o = 32'h05a68fd5 ;
			32'h00100288 : data_o = 32'h001006b7 ;
			32'h0010028c : data_o = 32'h8fcd8df5 ;
			32'h00100290 : data_o = 32'h06f7e793 ;
			32'h00100294 : data_o = 32'h100fc31c ;
			32'h00100298 : data_o = 32'h45010000 ;
			32'h0010029c : data_o = 32'h45058082 ;
			32'h001002a0 : data_o = 32'h20738082 ;
			32'h001002a4 : data_o = 32'h80823045 ;
			32'h001002a8 : data_o = 32'h30453073 ;
			32'h001002ac : data_o = 32'hc5098082 ;
			32'h001002b0 : data_o = 32'ha07347a1 ;
			32'h001002b4 : data_o = 32'h80823007 ;
			32'h001002b8 : data_o = 32'hb07347a1 ;
			32'h001002bc : data_o = 32'h80823007 ;
			32'h001002c0 : data_o = 32'hc6061141 ;
			32'h001002c4 : data_o = 32'h00000517 ;
			32'h001002c8 : data_o = 32'h31050513 ;
			32'h001002cc : data_o = 32'h05173dd5 ;
			32'h001002d0 : data_o = 32'h05130000 ;
			32'h001002d4 : data_o = 32'h35ed3165 ;
			32'h001002d8 : data_o = 32'h00000517 ;
			32'h001002dc : data_o = 32'h31c50513 ;
			32'h001002e0 : data_o = 32'h257335c5 ;
			32'h001002e4 : data_o = 32'h3df53410 ;
			32'h001002e8 : data_o = 32'h00000517 ;
			32'h001002ec : data_o = 32'h31850513 ;
			32'h001002f0 : data_o = 32'h25733dc1 ;
			32'h001002f4 : data_o = 32'h35f53420 ;
			32'h001002f8 : data_o = 32'h00000517 ;
			32'h001002fc : data_o = 32'h31450513 ;
			32'h00100300 : data_o = 32'h257335c1 ;
			32'h00100304 : data_o = 32'h3df13430 ;
			32'h00100308 : data_o = 32'h3db54529 ;
			32'h0010030c : data_o = 32'h1141a001 ;
			32'h00100310 : data_o = 32'h6541c606 ;
			32'h00100314 : data_o = 32'h45053779 ;
			32'h00100318 : data_o = 32'h40b23f59 ;
			32'h0010031c : data_o = 32'h80820141 ;
			32'h00100320 : data_o = 32'h8b85451c ;
			32'h00100324 : data_o = 32'h4108e399 ;
			32'h00100328 : data_o = 32'h557d8082 ;
			32'h0010032c : data_o = 32'h451c8082 ;
			32'h00100330 : data_o = 32'hfff58b89 ;
			32'h00100334 : data_o = 32'h8082c14c ;
			32'h00100338 : data_o = 32'h080027b7 ;
			32'h0010033c : data_o = 32'hc798577d ;
			32'h00100340 : data_o = 32'hc788c7cc ;
			32'h00100344 : data_o = 32'h80828082 ;
			32'h00100348 : data_o = 32'h080027b7 ;
			32'h0010034c : data_o = 32'h438843cc ;
			32'h00100350 : data_o = 32'h1de343d8 ;
			32'h00100354 : data_o = 32'h8082feb7 ;
			32'h00100358 : data_o = 32'hc686715d ;
			32'h0010035c : data_o = 32'hc29ac496 ;
			32'h00100360 : data_o = 32'hde22c09e ;
			32'h00100364 : data_o = 32'hda2adc26 ;
			32'h00100368 : data_o = 32'hd632d82e ;
			32'h0010036c : data_o = 32'hd23ad436 ;
			32'h00100370 : data_o = 32'hce42d03e ;
			32'h00100374 : data_o = 32'hca72cc46 ;
			32'h00100378 : data_o = 32'hc67ac876 ;
			32'h0010037c : data_o = 32'h0797c47e ;
			32'h00100380 : data_o = 32'h87930010 ;
			32'h00100384 : data_o = 32'h4380c927 ;
			32'h00100388 : data_o = 32'h3f7d43c4 ;
			32'h0010038c : data_o = 32'h34339522 ;
			32'h00100390 : data_o = 32'h95a60085 ;
			32'h00100394 : data_o = 32'h374d95a2 ;
			32'h00100398 : data_o = 32'h00100597 ;
			32'h0010039c : data_o = 32'hc8058593 ;
			32'h001003a0 : data_o = 32'h41c44180 ;
			32'h001003a4 : data_o = 32'h00140513 ;
			32'h001003a8 : data_o = 32'h00853633 ;
			32'h001003ac : data_o = 32'h009607b3 ;
			32'h001003b0 : data_o = 32'hc1dcc188 ;
			32'h001003b4 : data_o = 32'h42a640b6 ;
			32'h001003b8 : data_o = 32'h43864316 ;
			32'h001003bc : data_o = 32'h54e25472 ;
			32'h001003c0 : data_o = 32'h55c25552 ;
			32'h001003c4 : data_o = 32'h56a25632 ;
			32'h001003c8 : data_o = 32'h57825712 ;
			32'h001003cc : data_o = 32'h48e24872 ;
			32'h001003d0 : data_o = 32'h4ec24e52 ;
			32'h001003d4 : data_o = 32'h4fa24f32 ;
			32'h001003d8 : data_o = 32'h00736161 ;
			32'h001003dc : data_o = 32'h07973020 ;
			32'h001003e0 : data_o = 32'h87930010 ;
			32'h001003e4 : data_o = 32'h4388c3a7 ;
			32'h001003e8 : data_o = 32'h808243cc ;
			32'h001003ec : data_o = 32'hc6061141 ;
			32'h001003f0 : data_o = 32'hc226c422 ;
			32'h001003f4 : data_o = 32'h84ae842a ;
			32'h001003f8 : data_o = 32'h00100797 ;
			32'h001003fc : data_o = 32'hc2078793 ;
			32'h00100400 : data_o = 32'h47014681 ;
			32'h00100404 : data_o = 32'hc3d8c394 ;
			32'h00100408 : data_o = 32'h00100797 ;
			32'h0010040c : data_o = 32'hc0878793 ;
			32'h00100410 : data_o = 32'hc3ccc388 ;
			32'h00100414 : data_o = 32'h95223f15 ;
			32'h00100418 : data_o = 32'h00853433 ;
			32'h0010041c : data_o = 32'h95a295a6 ;
			32'h00100420 : data_o = 32'h05133f21 ;
			32'h00100424 : data_o = 32'h3db50800 ;
			32'h00100428 : data_o = 32'h35514505 ;
			32'h0010042c : data_o = 32'h442240b2 ;
			32'h00100430 : data_o = 32'h01414492 ;
			32'h00100434 : data_o = 32'h07938082 ;
			32'h00100438 : data_o = 32'hb0730800 ;
			32'h0010043c : data_o = 32'h80823047 ;
			32'h00100440 : data_o = 32'h8082c10c ;
			32'h00100444 : data_o = 32'h80824108 ;
			32'h00100448 : data_o = 32'h47854118 ;
			32'h0010044c : data_o = 32'h00b797b3 ;
			32'h00100450 : data_o = 32'hfff7c793 ;
			32'h00100454 : data_o = 32'h16338ff9 ;
			32'h00100458 : data_o = 32'h8e5d00b6 ;
			32'h0010045c : data_o = 32'h8082c110 ;
			32'h00100460 : data_o = 32'h55334108 ;
			32'h00100464 : data_o = 32'h890500b5 ;
			32'h00100468 : data_o = 32'h07b78082 ;
			32'h0010046c : data_o = 32'hcb887000 ;
			32'h00100470 : data_o = 32'h47838082 ;
			32'h00100474 : data_o = 32'h07a20015 ;
			32'h00100478 : data_o = 32'h00254703 ;
			32'h0010047c : data_o = 32'h8fd90742 ;
			32'h00100480 : data_o = 32'h00054703 ;
			32'h00100484 : data_o = 32'h47038fd9 ;
			32'h00100488 : data_o = 32'h07620035 ;
			32'h0010048c : data_o = 32'h07378fd9 ;
			32'h00100490 : data_o = 32'hcf1c7000 ;
			32'h00100494 : data_o = 32'h07b78082 ;
			32'h00100498 : data_o = 32'h47057000 ;
			32'h0010049c : data_o = 32'h8082d398 ;
			32'h001004a0 : data_o = 32'h70000737 ;
			32'h001004a4 : data_o = 32'hdffd535c ;
			32'h001004a8 : data_o = 32'h700007b7 ;
			32'h001004ac : data_o = 32'h80825788 ;
			32'h001004b0 : data_o = 32'hc6061141 ;
			32'h001004b4 : data_o = 32'h00020537 ;
			32'h001004b8 : data_o = 32'h450533ed ;
			32'h001004bc : data_o = 32'h07b73bcd ;
			32'h001004c0 : data_o = 32'h47057000 ;
			32'h001004c4 : data_o = 32'h40b2db98 ;
			32'h001004c8 : data_o = 32'h80820141 ;
			32'h001004cc : data_o = 32'hc6061141 ;
			32'h001004d0 : data_o = 32'h700007b7 ;
			32'h001004d4 : data_o = 32'h0207a823 ;
			32'h001004d8 : data_o = 32'h00020537 ;
			32'h001004dc : data_o = 32'h40b233f1 ;
			32'h001004e0 : data_o = 32'h80820141 ;
			32'h001004e4 : data_o = 32'h700007b7 ;
			32'h001004e8 : data_o = 32'h8082dbc8 ;
			32'h001004ec : data_o = 32'h00781141 ;
			32'h001004f0 : data_o = 32'h700007b7 ;
			32'h001004f4 : data_o = 32'h0141dfd8 ;
			32'h001004f8 : data_o = 32'h07b78082 ;
			32'h001004fc : data_o = 32'hdf887000 ;
			32'h00100500 : data_o = 32'h07b78082 ;
			32'h00100504 : data_o = 32'h43a87000 ;
			32'h00100508 : data_o = 32'h0ff57513 ;
			32'h0010050c : data_o = 32'h07b78082 ;
			32'h00100510 : data_o = 32'h47057000 ;
			32'h00100514 : data_o = 32'h8082c3f8 ;
			32'h00100518 : data_o = 32'h700007b7 ;
			32'h0010051c : data_o = 32'h0407a223 ;
			32'h00100520 : data_o = 32'h07b78082 ;
			32'h00100524 : data_o = 32'hc7a87000 ;
			32'h00100528 : data_o = 32'h07b78082 ;
			32'h0010052c : data_o = 32'hc7e87000 ;
			32'h00100530 : data_o = 32'h058e8082 ;
			32'h00100534 : data_o = 32'h8a1589e1 ;
			32'h00100538 : data_o = 32'h17b78dd1 ;
			32'h0010053c : data_o = 32'h87937000 ;
			32'h00100540 : data_o = 32'h8ddd8007 ;
			32'h00100544 : data_o = 32'hc793411c ;
			32'h00100548 : data_o = 32'hc19cfff7 ;
			32'h0010054c : data_o = 32'hf06f8082 ;
			32'h00100550 : data_o = 32'h0093d73f ;
			32'h00100554 : data_o = 32'h81060000 ;
			32'h00100558 : data_o = 32'h82068186 ;
			32'h0010055c : data_o = 32'h83068286 ;
			32'h00100560 : data_o = 32'h84068386 ;
			32'h00100564 : data_o = 32'h85068486 ;
			32'h00100568 : data_o = 32'h86068586 ;
			32'h0010056c : data_o = 32'h87068686 ;
			32'h00100570 : data_o = 32'h88068786 ;
			32'h00100574 : data_o = 32'h89068886 ;
			32'h00100578 : data_o = 32'h8a068986 ;
			32'h0010057c : data_o = 32'h8b068a86 ;
			32'h00100580 : data_o = 32'h8c068b86 ;
			32'h00100584 : data_o = 32'h8d068c86 ;
			32'h00100588 : data_o = 32'h8e068d86 ;
			32'h0010058c : data_o = 32'h8f068e86 ;
			32'h00100590 : data_o = 32'h01178f86 ;
			32'h00100594 : data_o = 32'h01130011 ;
			32'h00100598 : data_o = 32'h0d17a6e1 ;
			32'h0010059c : data_o = 32'h0d130010 ;
			32'h001005a0 : data_o = 32'h0d97a6ed ;
			32'h001005a4 : data_o = 32'h8d930010 ;
			32'h001005a8 : data_o = 32'h5763a7ed ;
			32'h001005ac : data_o = 32'h202301bd ;
			32'h001005b0 : data_o = 32'h0d11000d ;
			32'h001005b4 : data_o = 32'hffaddde3 ;
			32'h001005b8 : data_o = 32'h45814501 ;
			32'h001005bc : data_o = 32'hb75ff0ef ;
			32'h001005c0 : data_o = 32'h000202b7 ;
			32'h001005c4 : data_o = 32'h430502a1 ;
			32'h001005c8 : data_o = 32'h0062a023 ;
			32'h001005cc : data_o = 32'h10500073 ;
			32'h001005d0 : data_o = 32'h0000bff5 ;
			32'h001005d4 : data_o = 32'h45435845 ;
			32'h001005d8 : data_o = 32'h4f495450 ;
			32'h001005dc : data_o = 32'h2121214e ;
			32'h001005e0 : data_o = 32'h0000000a ;
			32'h001005e4 : data_o = 32'h3d3d3d3d ;
			32'h001005e8 : data_o = 32'h3d3d3d3d ;
			32'h001005ec : data_o = 32'h3d3d3d3d ;
			32'h001005f0 : data_o = 32'h0000000a ;
			32'h001005f4 : data_o = 32'h4350454d ;
			32'h001005f8 : data_o = 32'h2020203a ;
			32'h001005fc : data_o = 32'h00007830 ;
			32'h00100600 : data_o = 32'h41434d0a ;
			32'h00100604 : data_o = 32'h3a455355 ;
			32'h00100608 : data_o = 32'h00783020 ;
			32'h0010060c : data_o = 32'h56544d0a ;
			32'h00100610 : data_o = 32'h203a4c41 ;
			32'h00100614 : data_o = 32'h00783020 ;
			32'h00100618 : data_o = 32'h00100000 ;
			default : data_o = 32'h00000000 ;
		endcase 
	end
endmodule
