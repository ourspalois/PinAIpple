module rom_1p #(
	int Depth, 
 	int DATA_WIDTH = 32, 
 	int ADDR_WIDTH = 32 
 ) (
	input logic clk_i, 
	input logic req_i, 
	input logic [ADDR_WIDTH-1:0] addr_i, 
	output logic [DATA_WIDTH-1:0] data_o 
 );
	always_ff @(posedge clk_i) begin
		case (addr_i)
			32'h00100000 : data_o = 32'h3290006f ;
			32'h00100004 : data_o = 32'h3250006f ;
			32'h00100008 : data_o = 32'h3210006f ;
			32'h0010000c : data_o = 32'h31d0006f ;
			32'h00100010 : data_o = 32'h3190006f ;
			32'h00100014 : data_o = 32'h3150006f ;
			32'h00100018 : data_o = 32'h3110006f ;
			32'h0010001c : data_o = 32'h30d0006f ;
			32'h00100020 : data_o = 32'h3090006f ;
			32'h00100024 : data_o = 32'h3050006f ;
			32'h00100028 : data_o = 32'h3010006f ;
			32'h0010002c : data_o = 32'h2fd0006f ;
			32'h00100030 : data_o = 32'h2f90006f ;
			32'h00100034 : data_o = 32'h2f50006f ;
			32'h00100038 : data_o = 32'h2f10006f ;
			32'h0010003c : data_o = 32'h2ed0006f ;
			32'h00100040 : data_o = 32'h2e90006f ;
			32'h00100044 : data_o = 32'h0400006f ;
			32'h00100048 : data_o = 32'h2e10006f ;
			32'h0010004c : data_o = 32'h2dd0006f ;
			32'h00100050 : data_o = 32'h2d90006f ;
			32'h00100054 : data_o = 32'h2d50006f ;
			32'h00100058 : data_o = 32'h2d10006f ;
			32'h0010005c : data_o = 32'h2cd0006f ;
			32'h00100060 : data_o = 32'h2c90006f ;
			32'h00100064 : data_o = 32'h2c50006f ;
			32'h00100068 : data_o = 32'h2c10006f ;
			32'h0010006c : data_o = 32'h2bd0006f ;
			32'h00100070 : data_o = 32'h2b90006f ;
			32'h00100074 : data_o = 32'h2b50006f ;
			32'h00100078 : data_o = 32'h2b10006f ;
			32'h0010007c : data_o = 32'h2ad0006f ;
			32'h00100080 : data_o = 32'h07e0106f ;
			32'h00100084 : data_o = 32'hc686715d ;
			32'h00100088 : data_o = 32'hc29ac496 ;
			32'h0010008c : data_o = 32'hde22c09e ;
			32'h00100090 : data_o = 32'hda2edc2a ;
			32'h00100094 : data_o = 32'hd636d832 ;
			32'h00100098 : data_o = 32'hd23ed43a ;
			32'h0010009c : data_o = 32'hce46d042 ;
			32'h001000a0 : data_o = 32'hca76cc72 ;
			32'h001000a4 : data_o = 32'hc67ec87a ;
			32'h001000a8 : data_o = 32'h00ef0880 ;
			32'h001000ac : data_o = 32'h872a7510 ;
			32'h001000b0 : data_o = 32'h00100797 ;
			32'h001000b4 : data_o = 32'hf6478793 ;
			32'h001000b8 : data_o = 32'h0797c398 ;
			32'h001000bc : data_o = 32'h87930010 ;
			32'h001000c0 : data_o = 32'h4705f5e7 ;
			32'h001000c4 : data_o = 32'h0001c398 ;
			32'h001000c8 : data_o = 32'h42a640b6 ;
			32'h001000cc : data_o = 32'h43864316 ;
			32'h001000d0 : data_o = 32'h55625472 ;
			32'h001000d4 : data_o = 32'h564255d2 ;
			32'h001000d8 : data_o = 32'h572256b2 ;
			32'h001000dc : data_o = 32'h58025792 ;
			32'h001000e0 : data_o = 32'h4e6248f2 ;
			32'h001000e4 : data_o = 32'h4f424ed2 ;
			32'h001000e8 : data_o = 32'h61614fb2 ;
			32'h001000ec : data_o = 32'h30200073 ;
			32'h001000f0 : data_o = 32'hd6067179 ;
			32'h001000f4 : data_o = 32'h1800d422 ;
			32'h001000f8 : data_o = 32'hfca42e23 ;
			32'h001000fc : data_o = 32'hfe042623 ;
			32'h00100100 : data_o = 32'h2783a005 ;
			32'h00100104 : data_o = 32'h2703fec4 ;
			32'h00100108 : data_o = 32'h97bafdc4 ;
			32'h0010010c : data_o = 32'h0007c783 ;
			32'h00100110 : data_o = 32'h00ef853e ;
			32'h00100114 : data_o = 32'h27837640 ;
			32'h00100118 : data_o = 32'h0785fec4 ;
			32'h0010011c : data_o = 32'hfef42623 ;
			32'h00100120 : data_o = 32'hfec42783 ;
			32'h00100124 : data_o = 32'hfdc42703 ;
			32'h00100128 : data_o = 32'hc78397ba ;
			32'h0010012c : data_o = 32'hfbf10007 ;
			32'h00100130 : data_o = 32'h00010001 ;
			32'h00100134 : data_o = 32'h542250b2 ;
			32'h00100138 : data_o = 32'h80826145 ;
			32'h0010013c : data_o = 32'hd6067179 ;
			32'h00100140 : data_o = 32'h1800d422 ;
			32'h00100144 : data_o = 32'h8e2e8eaa ;
			32'h00100148 : data_o = 32'h85368332 ;
			32'h0010014c : data_o = 32'h863e85ba ;
			32'h00100150 : data_o = 32'h874686c2 ;
			32'h00100154 : data_o = 32'h0fa387f6 ;
			32'h00100158 : data_o = 32'h87f2fcf4 ;
			32'h0010015c : data_o = 32'hfcf40f23 ;
			32'h00100160 : data_o = 32'h0ea3879a ;
			32'h00100164 : data_o = 32'h87aafcf4 ;
			32'h00100168 : data_o = 32'hfcf40e23 ;
			32'h0010016c : data_o = 32'h0da387ae ;
			32'h00100170 : data_o = 32'h87b2fcf4 ;
			32'h00100174 : data_o = 32'hfcf40d23 ;
			32'h00100178 : data_o = 32'h0ca387b6 ;
			32'h0010017c : data_o = 32'h87bafcf4 ;
			32'h00100180 : data_o = 32'hfcf40c23 ;
			32'h00100184 : data_o = 32'h00ef4505 ;
			32'h00100188 : data_o = 32'h47836df0 ;
			32'h0010018c : data_o = 32'h9713fdf4 ;
			32'h00100190 : data_o = 32'h47830187 ;
			32'h00100194 : data_o = 32'h07c2fde4 ;
			32'h00100198 : data_o = 32'h47838f5d ;
			32'h0010019c : data_o = 32'h07a2fdd4 ;
			32'h001001a0 : data_o = 32'h47838f5d ;
			32'h001001a4 : data_o = 32'h8fd9fdc4 ;
			32'h001001a8 : data_o = 32'hfef42623 ;
			32'h001001ac : data_o = 32'hfd844783 ;
			32'h001001b0 : data_o = 32'h00ef853e ;
			32'h001001b4 : data_o = 32'h46836d10 ;
			32'h001001b8 : data_o = 32'h4703fd94 ;
			32'h001001bc : data_o = 32'h4783fda4 ;
			32'h001001c0 : data_o = 32'h863afdb4 ;
			32'h001001c4 : data_o = 32'h250385be ;
			32'h001001c8 : data_o = 32'h00effec4 ;
			32'h001001cc : data_o = 32'h00016d90 ;
			32'h001001d0 : data_o = 32'h542250b2 ;
			32'h001001d4 : data_o = 32'h80826145 ;
			32'h001001d8 : data_o = 32'hce061101 ;
			32'h001001dc : data_o = 32'h1000cc22 ;
			32'h001001e0 : data_o = 32'h8e2e8eaa ;
			32'h001001e4 : data_o = 32'h85368332 ;
			32'h001001e8 : data_o = 32'h863e85ba ;
			32'h001001ec : data_o = 32'h874686c2 ;
			32'h001001f0 : data_o = 32'h07a387f6 ;
			32'h001001f4 : data_o = 32'h87f2fef4 ;
			32'h001001f8 : data_o = 32'hfef40723 ;
			32'h001001fc : data_o = 32'h06a3879a ;
			32'h00100200 : data_o = 32'h87aafef4 ;
			32'h00100204 : data_o = 32'hfef40623 ;
			32'h00100208 : data_o = 32'h05a387ae ;
			32'h0010020c : data_o = 32'h87b2fef4 ;
			32'h00100210 : data_o = 32'hfef40523 ;
			32'h00100214 : data_o = 32'h04a387b6 ;
			32'h00100218 : data_o = 32'h87bafef4 ;
			32'h0010021c : data_o = 32'hfef40423 ;
			32'h00100220 : data_o = 32'h00ef4505 ;
			32'h00100224 : data_o = 32'h46834d50 ;
			32'h00100228 : data_o = 32'h4603fec4 ;
			32'h0010022c : data_o = 32'h4703fed4 ;
			32'h00100230 : data_o = 32'h4783fee4 ;
			32'h00100234 : data_o = 32'h85bafef4 ;
			32'h00100238 : data_o = 32'h00ef853e ;
			32'h0010023c : data_o = 32'h46834db0 ;
			32'h00100240 : data_o = 32'h4603fe84 ;
			32'h00100244 : data_o = 32'h4703fe94 ;
			32'h00100248 : data_o = 32'h4783fea4 ;
			32'h0010024c : data_o = 32'h85bafeb4 ;
			32'h00100250 : data_o = 32'h00ef853e ;
			32'h00100254 : data_o = 32'h401c5190 ;
			32'h00100258 : data_o = 32'h00ef853e ;
			32'h0010025c : data_o = 32'h00ef5670 ;
			32'h00100260 : data_o = 32'h401c5830 ;
			32'h00100264 : data_o = 32'h00efe789 ;
			32'h00100268 : data_o = 32'h87aa5950 ;
			32'h0010026c : data_o = 32'h4018a00d ;
			32'h00100270 : data_o = 32'h16634789 ;
			32'h00100274 : data_o = 32'h00ef00f7 ;
			32'h00100278 : data_o = 32'h87aa59d0 ;
			32'h0010027c : data_o = 32'h4018a809 ;
			32'h00100280 : data_o = 32'h16634785 ;
			32'h00100284 : data_o = 32'h00ef00f7 ;
			32'h00100288 : data_o = 32'h87aa5a50 ;
			32'h0010028c : data_o = 32'h853ea009 ;
			32'h00100290 : data_o = 32'h446240f2 ;
			32'h00100294 : data_o = 32'h80826105 ;
			32'h00100298 : data_o = 32'hd6067179 ;
			32'h0010029c : data_o = 32'h1800d422 ;
			32'h001002a0 : data_o = 32'h86ae87aa ;
			32'h001002a4 : data_o = 32'h0fa38732 ;
			32'h001002a8 : data_o = 32'h87b6fcf4 ;
			32'h001002ac : data_o = 32'hfcf40f23 ;
			32'h001002b0 : data_o = 32'h0ea387ba ;
			32'h001002b4 : data_o = 32'h4783fcf4 ;
			32'h001002b8 : data_o = 32'h078efdf4 ;
			32'h001002bc : data_o = 32'h0187f713 ;
			32'h001002c0 : data_o = 32'hfde44783 ;
			32'h001002c4 : data_o = 32'h8f5d0796 ;
			32'h001002c8 : data_o = 32'hfdd44783 ;
			32'h001002cc : data_o = 32'h8b91078a ;
			32'h001002d0 : data_o = 32'h26238fd9 ;
			32'h001002d4 : data_o = 32'h2503fef4 ;
			32'h001002d8 : data_o = 32'h00effec4 ;
			32'h001002dc : data_o = 32'h87aa5690 ;
			32'h001002e0 : data_o = 32'h50b2853e ;
			32'h001002e4 : data_o = 32'h61455422 ;
			32'h001002e8 : data_o = 32'h71798082 ;
			32'h001002ec : data_o = 32'hd422d606 ;
			32'h001002f0 : data_o = 32'h2e231800 ;
			32'h001002f4 : data_o = 32'h2783fca4 ;
			32'h001002f8 : data_o = 32'h2423fdc4 ;
			32'h001002fc : data_o = 32'h2623fef4 ;
			32'h00100300 : data_o = 32'ha835fe04 ;
			32'h00100304 : data_o = 32'hfe842703 ;
			32'h00100308 : data_o = 32'h77b347a9 ;
			32'h0010030c : data_o = 32'hf79302f7 ;
			32'h00100310 : data_o = 32'h87930ff7 ;
			32'h00100314 : data_o = 32'hf7130307 ;
			32'h00100318 : data_o = 32'h27830ff7 ;
			32'h0010031c : data_o = 32'h17c1fec4 ;
			32'h00100320 : data_o = 32'h8a2397a2 ;
			32'h00100324 : data_o = 32'h2703fee7 ;
			32'h00100328 : data_o = 32'h47a9fe84 ;
			32'h0010032c : data_o = 32'h02f757b3 ;
			32'h00100330 : data_o = 32'hfef42423 ;
			32'h00100334 : data_o = 32'hfec42783 ;
			32'h00100338 : data_o = 32'h26230785 ;
			32'h0010033c : data_o = 32'h2703fef4 ;
			32'h00100340 : data_o = 32'h478dfec4 ;
			32'h00100344 : data_o = 32'hfce7d0e3 ;
			32'h00100348 : data_o = 32'h2623478d ;
			32'h0010034c : data_o = 32'ha831fef4 ;
			32'h00100350 : data_o = 32'hfec42783 ;
			32'h00100354 : data_o = 32'h97a217c1 ;
			32'h00100358 : data_o = 32'hff47c783 ;
			32'h0010035c : data_o = 32'h2b21853e ;
			32'h00100360 : data_o = 32'hfec42783 ;
			32'h00100364 : data_o = 32'h262317fd ;
			32'h00100368 : data_o = 32'h2783fef4 ;
			32'h0010036c : data_o = 32'hd1e3fec4 ;
			32'h00100370 : data_o = 32'h0001fe07 ;
			32'h00100374 : data_o = 32'h50b20001 ;
			32'h00100378 : data_o = 32'h61455422 ;
			32'h0010037c : data_o = 32'h71798082 ;
			32'h00100380 : data_o = 32'h1800d622 ;
			32'h00100384 : data_o = 32'hfca42e23 ;
			32'h00100388 : data_o = 32'hfdc42703 ;
			32'h0010038c : data_o = 32'h06400793 ;
			32'h00100390 : data_o = 32'h02f707b3 ;
			32'h00100394 : data_o = 32'hfef42223 ;
			32'h00100398 : data_o = 32'hfe042423 ;
			32'h0010039c : data_o = 32'hfe042623 ;
			32'h001003a0 : data_o = 32'h2783a819 ;
			32'h001003a4 : data_o = 32'h0785fe84 ;
			32'h001003a8 : data_o = 32'hfef42423 ;
			32'h001003ac : data_o = 32'hfec42783 ;
			32'h001003b0 : data_o = 32'h26230785 ;
			32'h001003b4 : data_o = 32'h2703fef4 ;
			32'h001003b8 : data_o = 32'h2783fec4 ;
			32'h001003bc : data_o = 32'h62e3fe44 ;
			32'h001003c0 : data_o = 32'h2783fef7 ;
			32'h001003c4 : data_o = 32'h853efe84 ;
			32'h001003c8 : data_o = 32'h61455432 ;
			32'h001003cc : data_o = 32'h01138082 ;
			32'h001003d0 : data_o = 32'h2e23de01 ;
			32'h001003d4 : data_o = 32'h2c232011 ;
			32'h001003d8 : data_o = 32'h14002081 ;
			32'h001003dc : data_o = 32'h800007b7 ;
			32'h001003e0 : data_o = 32'hc3984705 ;
			32'h001003e4 : data_o = 32'h02000513 ;
			32'h001003e8 : data_o = 32'h05132179 ;
			32'h001003ec : data_o = 32'h21610740 ;
			32'h001003f0 : data_o = 32'h06500513 ;
			32'h001003f4 : data_o = 32'h05132149 ;
			32'h001003f8 : data_o = 32'h29b50730 ;
			32'h001003fc : data_o = 32'h07400513 ;
			32'h00100400 : data_o = 32'h4529299d ;
			32'h00100404 : data_o = 32'h1517298d ;
			32'h00100408 : data_o = 32'h05130000 ;
			32'h0010040c : data_o = 32'h31cdebe5 ;
			32'h00100410 : data_o = 32'h3e800513 ;
			32'h00100414 : data_o = 32'h262337ad ;
			32'h00100418 : data_o = 32'ha835fe04 ;
			32'h0010041c : data_o = 32'hfec42783 ;
			32'h00100420 : data_o = 32'h0ff7f793 ;
			32'h00100424 : data_o = 32'h48014885 ;
			32'h00100428 : data_o = 32'h46814701 ;
			32'h0010042c : data_o = 32'h45814601 ;
			32'h00100430 : data_o = 32'h33294501 ;
			32'h00100434 : data_o = 32'hfec42783 ;
			32'h00100438 : data_o = 32'h0ff7f793 ;
			32'h0010043c : data_o = 32'h48054885 ;
			32'h00100440 : data_o = 32'h46814701 ;
			32'h00100444 : data_o = 32'h45814601 ;
			32'h00100448 : data_o = 32'h39cd4501 ;
			32'h0010044c : data_o = 32'hfec42783 ;
			32'h00100450 : data_o = 32'h26230785 ;
			32'h00100454 : data_o = 32'h2703fef4 ;
			32'h00100458 : data_o = 32'h0793fec4 ;
			32'h0010045c : data_o = 32'hffe303f0 ;
			32'h00100460 : data_o = 32'h2623fae7 ;
			32'h00100464 : data_o = 32'ha0b1fe04 ;
			32'h00100468 : data_o = 32'hfec42783 ;
			32'h0010046c : data_o = 32'h0ff7f793 ;
			32'h00100470 : data_o = 32'h48014885 ;
			32'h00100474 : data_o = 32'h06934701 ;
			32'h00100478 : data_o = 32'h06130ff0 ;
			32'h0010047c : data_o = 32'h05930ff0 ;
			32'h00100480 : data_o = 32'h05130ff0 ;
			32'h00100484 : data_o = 32'h395d0ff0 ;
			32'h00100488 : data_o = 32'hfec42783 ;
			32'h0010048c : data_o = 32'h0ff7f793 ;
			32'h00100490 : data_o = 32'h48054885 ;
			32'h00100494 : data_o = 32'h06934701 ;
			32'h00100498 : data_o = 32'h06130ff0 ;
			32'h0010049c : data_o = 32'h05930ff0 ;
			32'h001004a0 : data_o = 32'h05130ff0 ;
			32'h001004a4 : data_o = 32'h39590ff0 ;
			32'h001004a8 : data_o = 32'hfec42783 ;
			32'h001004ac : data_o = 32'h26230785 ;
			32'h001004b0 : data_o = 32'h2703fef4 ;
			32'h001004b4 : data_o = 32'h0793fec4 ;
			32'h001004b8 : data_o = 32'hf7e303f0 ;
			32'h001004bc : data_o = 32'h1717fae7 ;
			32'h001004c0 : data_o = 32'h07130000 ;
			32'h001004c4 : data_o = 32'h0793e667 ;
			32'h001004c8 : data_o = 32'h86bade84 ;
			32'h001004cc : data_o = 32'h20000713 ;
			32'h001004d0 : data_o = 32'h85b6863a ;
			32'h001004d4 : data_o = 32'h00ef853e ;
			32'h001004d8 : data_o = 32'h15174a90 ;
			32'h001004dc : data_o = 32'h05130000 ;
			32'h001004e0 : data_o = 32'h3139dfa5 ;
			32'h001004e4 : data_o = 32'h3e800513 ;
			32'h001004e8 : data_o = 32'h24233d59 ;
			32'h001004ec : data_o = 32'ha871fe04 ;
			32'h001004f0 : data_o = 32'hfe842783 ;
			32'h001004f4 : data_o = 32'h17c1078e ;
			32'h001004f8 : data_o = 32'hc50397a2 ;
			32'h001004fc : data_o = 32'h2783df87 ;
			32'h00100500 : data_o = 32'h078efe84 ;
			32'h00100504 : data_o = 32'h97a217c1 ;
			32'h00100508 : data_o = 32'hdf97c583 ;
			32'h0010050c : data_o = 32'hfe842783 ;
			32'h00100510 : data_o = 32'h17c1078e ;
			32'h00100514 : data_o = 32'hc60397a2 ;
			32'h00100518 : data_o = 32'h2783dfa7 ;
			32'h0010051c : data_o = 32'h078efe84 ;
			32'h00100520 : data_o = 32'h97a217c1 ;
			32'h00100524 : data_o = 32'hdfb7c683 ;
			32'h00100528 : data_o = 32'hfe842783 ;
			32'h0010052c : data_o = 32'h0ff7f793 ;
			32'h00100530 : data_o = 32'h48014885 ;
			32'h00100534 : data_o = 32'h31194701 ;
			32'h00100538 : data_o = 32'hfe842783 ;
			32'h0010053c : data_o = 32'h17c1078e ;
			32'h00100540 : data_o = 32'hc50397a2 ;
			32'h00100544 : data_o = 32'h2783dfc7 ;
			32'h00100548 : data_o = 32'h078efe84 ;
			32'h0010054c : data_o = 32'h97a217c1 ;
			32'h00100550 : data_o = 32'hdfd7c583 ;
			32'h00100554 : data_o = 32'hfe842783 ;
			32'h00100558 : data_o = 32'h17c1078e ;
			32'h0010055c : data_o = 32'hc60397a2 ;
			32'h00100560 : data_o = 32'h2783dfe7 ;
			32'h00100564 : data_o = 32'h078efe84 ;
			32'h00100568 : data_o = 32'h97a217c1 ;
			32'h0010056c : data_o = 32'hdff7c683 ;
			32'h00100570 : data_o = 32'hfe842783 ;
			32'h00100574 : data_o = 32'h0ff7f793 ;
			32'h00100578 : data_o = 32'h48054885 ;
			32'h0010057c : data_o = 32'h3e7d4701 ;
			32'h00100580 : data_o = 32'hfe842783 ;
			32'h00100584 : data_o = 32'h24230785 ;
			32'h00100588 : data_o = 32'h2703fef4 ;
			32'h0010058c : data_o = 32'h0793fe84 ;
			32'h00100590 : data_o = 32'hffe303f0 ;
			32'h00100594 : data_o = 32'h1517f4e7 ;
			32'h00100598 : data_o = 32'h05130000 ;
			32'h0010059c : data_o = 32'h3e89d4a5 ;
			32'h001005a0 : data_o = 32'h3e800513 ;
			32'h001005a4 : data_o = 32'h24233be9 ;
			32'h001005a8 : data_o = 32'ha871fe04 ;
			32'h001005ac : data_o = 32'hfe842783 ;
			32'h001005b0 : data_o = 32'h17c1078e ;
			32'h001005b4 : data_o = 32'hc50397a2 ;
			32'h001005b8 : data_o = 32'h2783df87 ;
			32'h001005bc : data_o = 32'h078efe84 ;
			32'h001005c0 : data_o = 32'h97a217c1 ;
			32'h001005c4 : data_o = 32'hdf97c583 ;
			32'h001005c8 : data_o = 32'hfe842783 ;
			32'h001005cc : data_o = 32'h17c1078e ;
			32'h001005d0 : data_o = 32'hc60397a2 ;
			32'h001005d4 : data_o = 32'h2783dfa7 ;
			32'h001005d8 : data_o = 32'h078efe84 ;
			32'h001005dc : data_o = 32'h97a217c1 ;
			32'h001005e0 : data_o = 32'hdfb7c683 ;
			32'h001005e4 : data_o = 32'hfe842783 ;
			32'h001005e8 : data_o = 32'h0ff7f793 ;
			32'h001005ec : data_o = 32'h48014881 ;
			32'h001005f0 : data_o = 32'h36a94701 ;
			32'h001005f4 : data_o = 32'hfe842783 ;
			32'h001005f8 : data_o = 32'h17c1078e ;
			32'h001005fc : data_o = 32'hc50397a2 ;
			32'h00100600 : data_o = 32'h2783dfc7 ;
			32'h00100604 : data_o = 32'h078efe84 ;
			32'h00100608 : data_o = 32'h97a217c1 ;
			32'h0010060c : data_o = 32'hdfd7c583 ;
			32'h00100610 : data_o = 32'hfe842783 ;
			32'h00100614 : data_o = 32'h17c1078e ;
			32'h00100618 : data_o = 32'hc60397a2 ;
			32'h0010061c : data_o = 32'h2783dfe7 ;
			32'h00100620 : data_o = 32'h078efe84 ;
			32'h00100624 : data_o = 32'h97a217c1 ;
			32'h00100628 : data_o = 32'hdff7c683 ;
			32'h0010062c : data_o = 32'hfe842783 ;
			32'h00100630 : data_o = 32'h0ff7f793 ;
			32'h00100634 : data_o = 32'h48054881 ;
			32'h00100638 : data_o = 32'h36094701 ;
			32'h0010063c : data_o = 32'hfe842783 ;
			32'h00100640 : data_o = 32'h24230785 ;
			32'h00100644 : data_o = 32'h2703fef4 ;
			32'h00100648 : data_o = 32'h0793fe84 ;
			32'h0010064c : data_o = 32'hffe303f0 ;
			32'h00100650 : data_o = 32'h1517f4e7 ;
			32'h00100654 : data_o = 32'h05130000 ;
			32'h00100658 : data_o = 32'h3c59c9e5 ;
			32'h0010065c : data_o = 32'h3e800513 ;
			32'h00100660 : data_o = 32'h45293b39 ;
			32'h00100664 : data_o = 32'h15172c09 ;
			32'h00100668 : data_o = 32'h05130000 ;
			32'h0010066c : data_o = 32'h3449c9a5 ;
			32'h00100670 : data_o = 32'h15172a6d ;
			32'h00100674 : data_o = 32'h05130000 ;
			32'h00100678 : data_o = 32'h3c9dc9e5 ;
			32'h0010067c : data_o = 32'h800007b7 ;
			32'h00100680 : data_o = 32'hc3984709 ;
			32'h00100684 : data_o = 32'h00001517 ;
			32'h00100688 : data_o = 32'hc9850513 ;
			32'h0010068c : data_o = 32'h47813495 ;
			32'h00100690 : data_o = 32'h2083853e ;
			32'h00100694 : data_o = 32'h240321c1 ;
			32'h00100698 : data_o = 32'h01132181 ;
			32'h0010069c : data_o = 32'h80822201 ;
			32'h001006a0 : data_o = 32'hd6067179 ;
			32'h001006a4 : data_o = 32'h1800d422 ;
			32'h001006a8 : data_o = 32'h0fa387aa ;
			32'h001006ac : data_o = 32'h4783fcf4 ;
			32'h001006b0 : data_o = 32'h05a3fdf4 ;
			32'h001006b4 : data_o = 32'h2623fef4 ;
			32'h001006b8 : data_o = 32'ha835fe04 ;
			32'h001006bc : data_o = 32'hfeb44703 ;
			32'h001006c0 : data_o = 32'h77b347a9 ;
			32'h001006c4 : data_o = 32'hf79302f7 ;
			32'h001006c8 : data_o = 32'h87930ff7 ;
			32'h001006cc : data_o = 32'hf7130307 ;
			32'h001006d0 : data_o = 32'h27830ff7 ;
			32'h001006d4 : data_o = 32'h17c1fec4 ;
			32'h001006d8 : data_o = 32'h8a2397a2 ;
			32'h001006dc : data_o = 32'h4703fee7 ;
			32'h001006e0 : data_o = 32'h47a9feb4 ;
			32'h001006e4 : data_o = 32'h02f757b3 ;
			32'h001006e8 : data_o = 32'hfef405a3 ;
			32'h001006ec : data_o = 32'hfec42783 ;
			32'h001006f0 : data_o = 32'h26230785 ;
			32'h001006f4 : data_o = 32'h2703fef4 ;
			32'h001006f8 : data_o = 32'h478dfec4 ;
			32'h001006fc : data_o = 32'hfce7d0e3 ;
			32'h00100700 : data_o = 32'h2623478d ;
			32'h00100704 : data_o = 32'ha831fef4 ;
			32'h00100708 : data_o = 32'hfec42783 ;
			32'h0010070c : data_o = 32'h97a217c1 ;
			32'h00100710 : data_o = 32'hff47c783 ;
			32'h00100714 : data_o = 32'h2285853e ;
			32'h00100718 : data_o = 32'hfec42783 ;
			32'h0010071c : data_o = 32'h262317fd ;
			32'h00100720 : data_o = 32'h2783fef4 ;
			32'h00100724 : data_o = 32'hd1e3fec4 ;
			32'h00100728 : data_o = 32'h0001fe07 ;
			32'h0010072c : data_o = 32'h50b20001 ;
			32'h00100730 : data_o = 32'h61455422 ;
			32'h00100734 : data_o = 32'h715d8082 ;
			32'h00100738 : data_o = 32'hc4a2c686 ;
			32'h0010073c : data_o = 32'h0880c2a6 ;
			32'h00100740 : data_o = 32'hfaa42e23 ;
			32'h00100744 : data_o = 32'hfe0407a3 ;
			32'h00100748 : data_o = 32'h4783a881 ;
			32'h0010074c : data_o = 32'h8385fef4 ;
			32'h00100750 : data_o = 32'h0ff7f693 ;
			32'h00100754 : data_o = 32'hfbc42783 ;
			32'h00100758 : data_o = 32'h0ff7f593 ;
			32'h0010075c : data_o = 32'hfef44783 ;
			32'h00100760 : data_o = 32'h00178713 ;
			32'h00100764 : data_o = 32'h41f75793 ;
			32'h00100768 : data_o = 32'h973e83fd ;
			32'h0010076c : data_o = 32'h07b38b05 ;
			32'h00100770 : data_o = 32'hf79340f7 ;
			32'h00100774 : data_o = 32'h44830ff7 ;
			32'h00100778 : data_o = 32'h863efef4 ;
			32'h0010077c : data_o = 32'h3e298536 ;
			32'h00100780 : data_o = 32'h9793872a ;
			32'h00100784 : data_o = 32'h17c10024 ;
			32'h00100788 : data_o = 32'hac2397a2 ;
			32'h0010078c : data_o = 32'h4783fce7 ;
			32'h00100790 : data_o = 32'h0785fef4 ;
			32'h00100794 : data_o = 32'hfef407a3 ;
			32'h00100798 : data_o = 32'hfef44703 ;
			32'h0010079c : data_o = 32'hf6e3479d ;
			32'h001007a0 : data_o = 32'h07a3fae7 ;
			32'h001007a4 : data_o = 32'ha095fe04 ;
			32'h001007a8 : data_o = 32'hfef44783 ;
			32'h001007ac : data_o = 32'hf7938b85 ;
			32'h001007b0 : data_o = 32'he7990ff7 ;
			32'h001007b4 : data_o = 32'h02000513 ;
			32'h001007b8 : data_o = 32'h0513287d ;
			32'h001007bc : data_o = 32'h286507c0 ;
			32'h001007c0 : data_o = 32'h2423478d ;
			32'h001007c4 : data_o = 32'ha80dfef4 ;
			32'h001007c8 : data_o = 32'hfef44783 ;
			32'h001007cc : data_o = 32'h17c1078a ;
			32'h001007d0 : data_o = 32'ha70397a2 ;
			32'h001007d4 : data_o = 32'h2783fd87 ;
			32'h001007d8 : data_o = 32'h078efe84 ;
			32'h001007dc : data_o = 32'h00f757b3 ;
			32'h001007e0 : data_o = 32'h0ff7f793 ;
			32'h001007e4 : data_o = 32'h3d6d853e ;
			32'h001007e8 : data_o = 32'h07c00513 ;
			32'h001007ec : data_o = 32'h27832069 ;
			32'h001007f0 : data_o = 32'h17fdfe84 ;
			32'h001007f4 : data_o = 32'hfef42423 ;
			32'h001007f8 : data_o = 32'hfe842783 ;
			32'h001007fc : data_o = 32'hfc07d6e3 ;
			32'h00100800 : data_o = 32'hfef44783 ;
			32'h00100804 : data_o = 32'h07a30785 ;
			32'h00100808 : data_o = 32'h4703fef4 ;
			32'h0010080c : data_o = 32'h479dfef4 ;
			32'h00100810 : data_o = 32'hf8e7fce3 ;
			32'h00100814 : data_o = 32'h02000513 ;
			32'h00100818 : data_o = 32'h452928b9 ;
			32'h0010081c : data_o = 32'h000128a9 ;
			32'h00100820 : data_o = 32'h442640b6 ;
			32'h00100824 : data_o = 32'h61614496 ;
			32'h00100828 : data_o = 32'h11018082 ;
			32'h0010082c : data_o = 32'hcc22ce06 ;
			32'h00100830 : data_o = 32'h26231000 ;
			32'h00100834 : data_o = 32'ha025fe04 ;
			32'h00100838 : data_o = 32'hfec42783 ;
			32'h0010083c : data_o = 32'h03f7f793 ;
			32'h00100840 : data_o = 32'h2783e791 ;
			32'h00100844 : data_o = 32'hc399fec4 ;
			32'h00100848 : data_o = 32'h20354529 ;
			32'h0010084c : data_o = 32'hfec42783 ;
			32'h00100850 : data_o = 32'h35d5853e ;
			32'h00100854 : data_o = 32'hfec42783 ;
			32'h00100858 : data_o = 32'h26230785 ;
			32'h0010085c : data_o = 32'h2703fef4 ;
			32'h00100860 : data_o = 32'h0793fec4 ;
			32'h00100864 : data_o = 32'hd9e30ff0 ;
			32'h00100868 : data_o = 32'h0001fce7 ;
			32'h0010086c : data_o = 32'h40f20001 ;
			32'h00100870 : data_o = 32'h61054462 ;
			32'h00100874 : data_o = 32'h11018082 ;
			32'h00100878 : data_o = 32'hcc22ce06 ;
			32'h0010087c : data_o = 32'h87aa1000 ;
			32'h00100880 : data_o = 32'hfef407a3 ;
			32'h00100884 : data_o = 32'hfef44703 ;
			32'h00100888 : data_o = 32'h166347a9 ;
			32'h0010088c : data_o = 32'h45b500f7 ;
			32'h00100890 : data_o = 32'h80001537 ;
			32'h00100894 : data_o = 32'h47832e2d ;
			32'h00100898 : data_o = 32'h85befef4 ;
			32'h0010089c : data_o = 32'h80001537 ;
			32'h001008a0 : data_o = 32'h4783263d ;
			32'h001008a4 : data_o = 32'h853efef4 ;
			32'h001008a8 : data_o = 32'h446240f2 ;
			32'h001008ac : data_o = 32'h80826105 ;
			32'h001008b0 : data_o = 32'hc6061141 ;
			32'h001008b4 : data_o = 32'h0800c422 ;
			32'h001008b8 : data_o = 32'h80001537 ;
			32'h001008bc : data_o = 32'h87aa24c5 ;
			32'h001008c0 : data_o = 32'h40b2853e ;
			32'h001008c4 : data_o = 32'h01414422 ;
			32'h001008c8 : data_o = 32'h11018082 ;
			32'h001008cc : data_o = 32'hcc22ce06 ;
			32'h001008d0 : data_o = 32'h26231000 ;
			32'h001008d4 : data_o = 32'ha819fea4 ;
			32'h001008d8 : data_o = 32'hfec42783 ;
			32'h001008dc : data_o = 32'h00178713 ;
			32'h001008e0 : data_o = 32'hfee42623 ;
			32'h001008e4 : data_o = 32'h0007c783 ;
			32'h001008e8 : data_o = 32'h3771853e ;
			32'h001008ec : data_o = 32'hfec42783 ;
			32'h001008f0 : data_o = 32'h0007c783 ;
			32'h001008f4 : data_o = 32'h4781f3f5 ;
			32'h001008f8 : data_o = 32'h40f2853e ;
			32'h001008fc : data_o = 32'h61054462 ;
			32'h00100900 : data_o = 32'h71798082 ;
			32'h00100904 : data_o = 32'hd422d606 ;
			32'h00100908 : data_o = 32'h2e231800 ;
			32'h0010090c : data_o = 32'h2623fca4 ;
			32'h00100910 : data_o = 32'ha891fe04 ;
			32'h00100914 : data_o = 32'hfdc42783 ;
			32'h00100918 : data_o = 32'h242383f1 ;
			32'h0010091c : data_o = 32'h2703fef4 ;
			32'h00100920 : data_o = 32'h47a5fe84 ;
			32'h00100924 : data_o = 32'h00e7cd63 ;
			32'h00100928 : data_o = 32'hfe842783 ;
			32'h0010092c : data_o = 32'h0ff7f793 ;
			32'h00100930 : data_o = 32'h03078793 ;
			32'h00100934 : data_o = 32'h0ff7f793 ;
			32'h00100938 : data_o = 32'h3f35853e ;
			32'h0010093c : data_o = 32'h2783a819 ;
			32'h00100940 : data_o = 32'hf793fe84 ;
			32'h00100944 : data_o = 32'h87930ff7 ;
			32'h00100948 : data_o = 32'hf7930377 ;
			32'h0010094c : data_o = 32'h853e0ff7 ;
			32'h00100950 : data_o = 32'h2783371d ;
			32'h00100954 : data_o = 32'h0792fdc4 ;
			32'h00100958 : data_o = 32'hfcf42e23 ;
			32'h0010095c : data_o = 32'hfec42783 ;
			32'h00100960 : data_o = 32'h26230785 ;
			32'h00100964 : data_o = 32'h2703fef4 ;
			32'h00100968 : data_o = 32'h479dfec4 ;
			32'h0010096c : data_o = 32'hfae7d4e3 ;
			32'h00100970 : data_o = 32'h00010001 ;
			32'h00100974 : data_o = 32'h542250b2 ;
			32'h00100978 : data_o = 32'h80826145 ;
			32'h0010097c : data_o = 32'hc6221141 ;
			32'h00100980 : data_o = 32'h07b70800 ;
			32'h00100984 : data_o = 32'h07a10002 ;
			32'h00100988 : data_o = 32'hc3984705 ;
			32'h0010098c : data_o = 32'h44320001 ;
			32'h00100990 : data_o = 32'h80820141 ;
			32'h00100994 : data_o = 32'hce221101 ;
			32'h00100998 : data_o = 32'h27f31000 ;
			32'h0010099c : data_o = 32'h26233410 ;
			32'h001009a0 : data_o = 32'h2783fef4 ;
			32'h001009a4 : data_o = 32'h853efec4 ;
			32'h001009a8 : data_o = 32'h61054472 ;
			32'h001009ac : data_o = 32'h11018082 ;
			32'h001009b0 : data_o = 32'h1000ce22 ;
			32'h001009b4 : data_o = 32'h342027f3 ;
			32'h001009b8 : data_o = 32'hfef42623 ;
			32'h001009bc : data_o = 32'hfec42783 ;
			32'h001009c0 : data_o = 32'h4472853e ;
			32'h001009c4 : data_o = 32'h80826105 ;
			32'h001009c8 : data_o = 32'hce221101 ;
			32'h001009cc : data_o = 32'h27f31000 ;
			32'h001009d0 : data_o = 32'h26233430 ;
			32'h001009d4 : data_o = 32'h2783fef4 ;
			32'h001009d8 : data_o = 32'h853efec4 ;
			32'h001009dc : data_o = 32'h61054472 ;
			32'h001009e0 : data_o = 32'h11018082 ;
			32'h001009e4 : data_o = 32'h1000ce22 ;
			32'h001009e8 : data_o = 32'hb00027f3 ;
			32'h001009ec : data_o = 32'hfef42623 ;
			32'h001009f0 : data_o = 32'hfec42783 ;
			32'h001009f4 : data_o = 32'h4472853e ;
			32'h001009f8 : data_o = 32'h80826105 ;
			32'h001009fc : data_o = 32'hc6221141 ;
			32'h00100a00 : data_o = 32'h10730800 ;
			32'h00100a04 : data_o = 32'h0001b000 ;
			32'h00100a08 : data_o = 32'h01414432 ;
			32'h00100a0c : data_o = 32'h71798082 ;
			32'h00100a10 : data_o = 32'h1800d622 ;
			32'h00100a14 : data_o = 32'hfca42e23 ;
			32'h00100a18 : data_o = 32'hfcb42c23 ;
			32'h00100a1c : data_o = 32'hfdc42703 ;
			32'h00100a20 : data_o = 32'hf46347fd ;
			32'h00100a24 : data_o = 32'h478500e7 ;
			32'h00100a28 : data_o = 32'hf797a879 ;
			32'h00100a2c : data_o = 32'h8793000f ;
			32'h00100a30 : data_o = 32'h43985d67 ;
			32'h00100a34 : data_o = 32'hfdc42783 ;
			32'h00100a38 : data_o = 32'h97ba078a ;
			32'h00100a3c : data_o = 32'hfef42623 ;
			32'h00100a40 : data_o = 32'hfd842703 ;
			32'h00100a44 : data_o = 32'hfec42783 ;
			32'h00100a48 : data_o = 32'h40f707b3 ;
			32'h00100a4c : data_o = 32'hfef42423 ;
			32'h00100a50 : data_o = 32'hfe842703 ;
			32'h00100a54 : data_o = 32'h000807b7 ;
			32'h00100a58 : data_o = 32'h00f75863 ;
			32'h00100a5c : data_o = 32'hfe842703 ;
			32'h00100a60 : data_o = 32'hfff807b7 ;
			32'h00100a64 : data_o = 32'h00f75463 ;
			32'h00100a68 : data_o = 32'ha8b14789 ;
			32'h00100a6c : data_o = 32'hfe842783 ;
			32'h00100a70 : data_o = 32'hfef42223 ;
			32'h00100a74 : data_o = 32'hfe442783 ;
			32'h00100a78 : data_o = 32'h01479713 ;
			32'h00100a7c : data_o = 32'h7fe007b7 ;
			32'h00100a80 : data_o = 32'h27838f7d ;
			32'h00100a84 : data_o = 32'h9693fe44 ;
			32'h00100a88 : data_o = 32'h07b70097 ;
			32'h00100a8c : data_o = 32'h8ff50010 ;
			32'h00100a90 : data_o = 32'h26838f5d ;
			32'h00100a94 : data_o = 32'hf7b7fe44 ;
			32'h00100a98 : data_o = 32'h8ff5000f ;
			32'h00100a9c : data_o = 32'h27838f5d ;
			32'h00100aa0 : data_o = 32'h9693fe44 ;
			32'h00100aa4 : data_o = 32'h07b700b7 ;
			32'h00100aa8 : data_o = 32'h8ff58000 ;
			32'h00100aac : data_o = 32'he7938fd9 ;
			32'h00100ab0 : data_o = 32'h202306f7 ;
			32'h00100ab4 : data_o = 32'h2783fef4 ;
			32'h00100ab8 : data_o = 32'h2703fec4 ;
			32'h00100abc : data_o = 32'hc398fe04 ;
			32'h00100ac0 : data_o = 32'h0000100f ;
			32'h00100ac4 : data_o = 32'h853e4781 ;
			32'h00100ac8 : data_o = 32'h61455432 ;
			32'h00100acc : data_o = 32'h11018082 ;
			32'h00100ad0 : data_o = 32'h1000ce22 ;
			32'h00100ad4 : data_o = 32'hfea42623 ;
			32'h00100ad8 : data_o = 32'hfec42783 ;
			32'h00100adc : data_o = 32'h3047a073 ;
			32'h00100ae0 : data_o = 32'h44720001 ;
			32'h00100ae4 : data_o = 32'h80826105 ;
			32'h00100ae8 : data_o = 32'hce221101 ;
			32'h00100aec : data_o = 32'h26231000 ;
			32'h00100af0 : data_o = 32'h2783fea4 ;
			32'h00100af4 : data_o = 32'hb073fec4 ;
			32'h00100af8 : data_o = 32'h00013047 ;
			32'h00100afc : data_o = 32'h61054472 ;
			32'h00100b00 : data_o = 32'h11018082 ;
			32'h00100b04 : data_o = 32'h1000ce22 ;
			32'h00100b08 : data_o = 32'hfea42623 ;
			32'h00100b0c : data_o = 32'hfec42783 ;
			32'h00100b10 : data_o = 32'h47a1c789 ;
			32'h00100b14 : data_o = 32'h3007a073 ;
			32'h00100b18 : data_o = 32'h47a1a021 ;
			32'h00100b1c : data_o = 32'h3007b073 ;
			32'h00100b20 : data_o = 32'h44720001 ;
			32'h00100b24 : data_o = 32'h80826105 ;
			32'h00100b28 : data_o = 32'hc6061141 ;
			32'h00100b2c : data_o = 32'h0800c422 ;
			32'h00100b30 : data_o = 32'h00001517 ;
			32'h00100b34 : data_o = 32'h9f450513 ;
			32'h00100b38 : data_o = 32'h15173b49 ;
			32'h00100b3c : data_o = 32'h05130000 ;
			32'h00100b40 : data_o = 32'h33619fa5 ;
			32'h00100b44 : data_o = 32'h00001517 ;
			32'h00100b48 : data_o = 32'ha0050513 ;
			32'h00100b4c : data_o = 32'h35993bbd ;
			32'h00100b50 : data_o = 32'h853e87aa ;
			32'h00100b54 : data_o = 32'h1517337d ;
			32'h00100b58 : data_o = 32'h05130000 ;
			32'h00100b5c : data_o = 32'h33b59fa5 ;
			32'h00100b60 : data_o = 32'h87aa35b9 ;
			32'h00100b64 : data_o = 32'h3b71853e ;
			32'h00100b68 : data_o = 32'h00001517 ;
			32'h00100b6c : data_o = 32'h9f450513 ;
			32'h00100b70 : data_o = 32'h3d993ba9 ;
			32'h00100b74 : data_o = 32'h853e87aa ;
			32'h00100b78 : data_o = 32'h45293369 ;
			32'h00100b7c : data_o = 32'h000139ed ;
			32'h00100b80 : data_o = 32'h1141bffd ;
			32'h00100b84 : data_o = 32'hc422c606 ;
			32'h00100b88 : data_o = 32'h65410800 ;
			32'h00100b8c : data_o = 32'h45053789 ;
			32'h00100b90 : data_o = 32'h00013f8d ;
			32'h00100b94 : data_o = 32'h442240b2 ;
			32'h00100b98 : data_o = 32'h80820141 ;
			32'h00100b9c : data_o = 32'hd6227179 ;
			32'h00100ba0 : data_o = 32'h2e231800 ;
			32'h00100ba4 : data_o = 32'h57fdfca4 ;
			32'h00100ba8 : data_o = 32'hfef42623 ;
			32'h00100bac : data_o = 32'hfdc42783 ;
			32'h00100bb0 : data_o = 32'h439c07a1 ;
			32'h00100bb4 : data_o = 32'he7918b85 ;
			32'h00100bb8 : data_o = 32'hfdc42783 ;
			32'h00100bbc : data_o = 32'h2623439c ;
			32'h00100bc0 : data_o = 32'h2783fef4 ;
			32'h00100bc4 : data_o = 32'h853efec4 ;
			32'h00100bc8 : data_o = 32'h61455432 ;
			32'h00100bcc : data_o = 32'h11018082 ;
			32'h00100bd0 : data_o = 32'h1000ce22 ;
			32'h00100bd4 : data_o = 32'hfea42623 ;
			32'h00100bd8 : data_o = 32'h05a387ae ;
			32'h00100bdc : data_o = 32'h0001fef4 ;
			32'h00100be0 : data_o = 32'hfec42783 ;
			32'h00100be4 : data_o = 32'h439c07a1 ;
			32'h00100be8 : data_o = 32'hfbfd8b89 ;
			32'h00100bec : data_o = 32'hfec42783 ;
			32'h00100bf0 : data_o = 32'h47030791 ;
			32'h00100bf4 : data_o = 32'hc398feb4 ;
			32'h00100bf8 : data_o = 32'h44720001 ;
			32'h00100bfc : data_o = 32'h80826105 ;
			32'h00100c00 : data_o = 32'hce221101 ;
			32'h00100c04 : data_o = 32'h24231000 ;
			32'h00100c08 : data_o = 32'h2623fea4 ;
			32'h00100c0c : data_o = 32'h26b7feb4 ;
			32'h00100c10 : data_o = 32'h06a10800 ;
			32'h00100c14 : data_o = 32'hc290567d ;
			32'h00100c18 : data_o = 32'hfec42683 ;
			32'h00100c1c : data_o = 32'h0006d713 ;
			32'h00100c20 : data_o = 32'h26b74781 ;
			32'h00100c24 : data_o = 32'h06b10800 ;
			32'h00100c28 : data_o = 32'hc29c87ba ;
			32'h00100c2c : data_o = 32'h080027b7 ;
			32'h00100c30 : data_o = 32'h270307a1 ;
			32'h00100c34 : data_o = 32'hc398fe84 ;
			32'h00100c38 : data_o = 32'h44720001 ;
			32'h00100c3c : data_o = 32'h80826105 ;
			32'h00100c40 : data_o = 32'hd6067179 ;
			32'h00100c44 : data_o = 32'h1800d422 ;
			32'h00100c48 : data_o = 32'hfca42c23 ;
			32'h00100c4c : data_o = 32'hfcb42e23 ;
			32'h00100c50 : data_o = 32'h242320fd ;
			32'h00100c54 : data_o = 32'h2623fea4 ;
			32'h00100c58 : data_o = 32'h2603feb4 ;
			32'h00100c5c : data_o = 32'h2683fe84 ;
			32'h00100c60 : data_o = 32'h2503fec4 ;
			32'h00100c64 : data_o = 32'h2583fd84 ;
			32'h00100c68 : data_o = 32'h0733fdc4 ;
			32'h00100c6c : data_o = 32'h883a00a6 ;
			32'h00100c70 : data_o = 32'h00c83833 ;
			32'h00100c74 : data_o = 32'h00b687b3 ;
			32'h00100c78 : data_o = 32'h00f806b3 ;
			32'h00100c7c : data_o = 32'h242387b6 ;
			32'h00100c80 : data_o = 32'h2623fee4 ;
			32'h00100c84 : data_o = 32'h2503fef4 ;
			32'h00100c88 : data_o = 32'h2583fe84 ;
			32'h00100c8c : data_o = 32'h3f8dfec4 ;
			32'h00100c90 : data_o = 32'h50b20001 ;
			32'h00100c94 : data_o = 32'h61455422 ;
			32'h00100c98 : data_o = 32'h715d8082 ;
			32'h00100c9c : data_o = 32'hc496c686 ;
			32'h00100ca0 : data_o = 32'hc09ec29a ;
			32'h00100ca4 : data_o = 32'hdc2ade22 ;
			32'h00100ca8 : data_o = 32'hd832da2e ;
			32'h00100cac : data_o = 32'hd43ad636 ;
			32'h00100cb0 : data_o = 32'hd042d23e ;
			32'h00100cb4 : data_o = 32'hcc72ce46 ;
			32'h00100cb8 : data_o = 32'hc87aca76 ;
			32'h00100cbc : data_o = 32'h0880c67e ;
			32'h00100cc0 : data_o = 32'h000ff797 ;
			32'h00100cc4 : data_o = 32'h36878793 ;
			32'h00100cc8 : data_o = 32'h43dc4398 ;
			32'h00100ccc : data_o = 32'h85be853a ;
			32'h00100cd0 : data_o = 32'hf7973f85 ;
			32'h00100cd4 : data_o = 32'h8793000f ;
			32'h00100cd8 : data_o = 32'h439834e7 ;
			32'h00100cdc : data_o = 32'h450543dc ;
			32'h00100ce0 : data_o = 32'h06334581 ;
			32'h00100ce4 : data_o = 32'h883200a7 ;
			32'h00100ce8 : data_o = 32'h00e83833 ;
			32'h00100cec : data_o = 32'h00b786b3 ;
			32'h00100cf0 : data_o = 32'h00d807b3 ;
			32'h00100cf4 : data_o = 32'h873286be ;
			32'h00100cf8 : data_o = 32'hf69787b6 ;
			32'h00100cfc : data_o = 32'h8693000f ;
			32'h00100d00 : data_o = 32'hc2983266 ;
			32'h00100d04 : data_o = 32'h0001c2dc ;
			32'h00100d08 : data_o = 32'h42a640b6 ;
			32'h00100d0c : data_o = 32'h43864316 ;
			32'h00100d10 : data_o = 32'h55625472 ;
			32'h00100d14 : data_o = 32'h564255d2 ;
			32'h00100d18 : data_o = 32'h572256b2 ;
			32'h00100d1c : data_o = 32'h58025792 ;
			32'h00100d20 : data_o = 32'h4e6248f2 ;
			32'h00100d24 : data_o = 32'h4f424ed2 ;
			32'h00100d28 : data_o = 32'h61614fb2 ;
			32'h00100d2c : data_o = 32'h30200073 ;
			32'h00100d30 : data_o = 32'hc6221141 ;
			32'h00100d34 : data_o = 32'h00010800 ;
			32'h00100d38 : data_o = 32'h01414432 ;
			32'h00100d3c : data_o = 32'h11018082 ;
			32'h00100d40 : data_o = 32'h1000ce22 ;
			32'h00100d44 : data_o = 32'h08002837 ;
			32'h00100d48 : data_o = 32'h28030811 ;
			32'h00100d4c : data_o = 32'h26230008 ;
			32'h00100d50 : data_o = 32'h2837ff04 ;
			32'h00100d54 : data_o = 32'h28030800 ;
			32'h00100d58 : data_o = 32'h24230008 ;
			32'h00100d5c : data_o = 32'h2837ff04 ;
			32'h00100d60 : data_o = 32'h08110800 ;
			32'h00100d64 : data_o = 32'h00082803 ;
			32'h00100d68 : data_o = 32'hfec42883 ;
			32'h00100d6c : data_o = 32'hfd089ce3 ;
			32'h00100d70 : data_o = 32'hfec42803 ;
			32'h00100d74 : data_o = 32'h45818542 ;
			32'h00100d78 : data_o = 32'h00051793 ;
			32'h00100d7c : data_o = 32'h25834701 ;
			32'h00100d80 : data_o = 32'h862efe84 ;
			32'h00100d84 : data_o = 32'h65b34681 ;
			32'h00100d88 : data_o = 32'h202300c7 ;
			32'h00100d8c : data_o = 32'h8fd5feb4 ;
			32'h00100d90 : data_o = 32'hfef42223 ;
			32'h00100d94 : data_o = 32'hfe042703 ;
			32'h00100d98 : data_o = 32'hfe442783 ;
			32'h00100d9c : data_o = 32'h85be853a ;
			32'h00100da0 : data_o = 32'h61054472 ;
			32'h00100da4 : data_o = 32'h11418082 ;
			32'h00100da8 : data_o = 32'h0800c622 ;
			32'h00100dac : data_o = 32'h000ff797 ;
			32'h00100db0 : data_o = 32'h27478793 ;
			32'h00100db4 : data_o = 32'h43dc4398 ;
			32'h00100db8 : data_o = 32'h85be853a ;
			32'h00100dbc : data_o = 32'h01414432 ;
			32'h00100dc0 : data_o = 32'h11018082 ;
			32'h00100dc4 : data_o = 32'hcc22ce06 ;
			32'h00100dc8 : data_o = 32'h24231000 ;
			32'h00100dcc : data_o = 32'h2623fea4 ;
			32'h00100dd0 : data_o = 32'hf797feb4 ;
			32'h00100dd4 : data_o = 32'h8793000f ;
			32'h00100dd8 : data_o = 32'h468124e7 ;
			32'h00100ddc : data_o = 32'hc3944701 ;
			32'h00100de0 : data_o = 32'hf697c3d8 ;
			32'h00100de4 : data_o = 32'h8693000f ;
			32'h00100de8 : data_o = 32'h27032466 ;
			32'h00100dec : data_o = 32'h2783fe84 ;
			32'h00100df0 : data_o = 32'hc298fec4 ;
			32'h00100df4 : data_o = 32'h2503c2dc ;
			32'h00100df8 : data_o = 32'h2583fe84 ;
			32'h00100dfc : data_o = 32'h3589fec4 ;
			32'h00100e00 : data_o = 32'h08000513 ;
			32'h00100e04 : data_o = 32'h450531e9 ;
			32'h00100e08 : data_o = 32'h000139ed ;
			32'h00100e0c : data_o = 32'h446240f2 ;
			32'h00100e10 : data_o = 32'h80826105 ;
			32'h00100e14 : data_o = 32'hc6221141 ;
			32'h00100e18 : data_o = 32'h07930800 ;
			32'h00100e1c : data_o = 32'hb0730800 ;
			32'h00100e20 : data_o = 32'h00013047 ;
			32'h00100e24 : data_o = 32'h01414432 ;
			32'h00100e28 : data_o = 32'h11018082 ;
			32'h00100e2c : data_o = 32'h1000ce22 ;
			32'h00100e30 : data_o = 32'hfea42623 ;
			32'h00100e34 : data_o = 32'hfeb42423 ;
			32'h00100e38 : data_o = 32'hfec42783 ;
			32'h00100e3c : data_o = 32'hfe842703 ;
			32'h00100e40 : data_o = 32'h0001c398 ;
			32'h00100e44 : data_o = 32'h61054472 ;
			32'h00100e48 : data_o = 32'h11018082 ;
			32'h00100e4c : data_o = 32'h1000ce22 ;
			32'h00100e50 : data_o = 32'hfea42623 ;
			32'h00100e54 : data_o = 32'hfec42783 ;
			32'h00100e58 : data_o = 32'h853e439c ;
			32'h00100e5c : data_o = 32'h61054472 ;
			32'h00100e60 : data_o = 32'h71798082 ;
			32'h00100e64 : data_o = 32'hd422d606 ;
			32'h00100e68 : data_o = 32'h2e231800 ;
			32'h00100e6c : data_o = 32'h2c23fca4 ;
			32'h00100e70 : data_o = 32'h2a23fcb4 ;
			32'h00100e74 : data_o = 32'h2503fcc4 ;
			32'h00100e78 : data_o = 32'h3fc1fdc4 ;
			32'h00100e7c : data_o = 32'hfea42623 ;
			32'h00100e80 : data_o = 32'hfd842783 ;
			32'h00100e84 : data_o = 32'h17b34705 ;
			32'h00100e88 : data_o = 32'hc79300f7 ;
			32'h00100e8c : data_o = 32'h873efff7 ;
			32'h00100e90 : data_o = 32'hfec42783 ;
			32'h00100e94 : data_o = 32'h26238ff9 ;
			32'h00100e98 : data_o = 32'h2783fef4 ;
			32'h00100e9c : data_o = 32'h2703fd84 ;
			32'h00100ea0 : data_o = 32'h17b3fd44 ;
			32'h00100ea4 : data_o = 32'h270300f7 ;
			32'h00100ea8 : data_o = 32'h8fd9fec4 ;
			32'h00100eac : data_o = 32'hfef42623 ;
			32'h00100eb0 : data_o = 32'hfec42583 ;
			32'h00100eb4 : data_o = 32'hfdc42503 ;
			32'h00100eb8 : data_o = 32'h00013f8d ;
			32'h00100ebc : data_o = 32'h542250b2 ;
			32'h00100ec0 : data_o = 32'h80826145 ;
			32'h00100ec4 : data_o = 32'hd6067179 ;
			32'h00100ec8 : data_o = 32'h1800d422 ;
			32'h00100ecc : data_o = 32'hfca42e23 ;
			32'h00100ed0 : data_o = 32'hfcb42c23 ;
			32'h00100ed4 : data_o = 32'hfdc42503 ;
			32'h00100ed8 : data_o = 32'h26233f8d ;
			32'h00100edc : data_o = 32'h2783fea4 ;
			32'h00100ee0 : data_o = 32'h2703fd84 ;
			32'h00100ee4 : data_o = 32'h57b3fec4 ;
			32'h00100ee8 : data_o = 32'h8b8500f7 ;
			32'h00100eec : data_o = 32'h50b2853e ;
			32'h00100ef0 : data_o = 32'h61455422 ;
			32'h00100ef4 : data_o = 32'h11018082 ;
			32'h00100ef8 : data_o = 32'h1000ce22 ;
			32'h00100efc : data_o = 32'hfea42623 ;
			32'h00100f00 : data_o = 32'h700007b7 ;
			32'h00100f04 : data_o = 32'h270307c1 ;
			32'h00100f08 : data_o = 32'hc398fec4 ;
			32'h00100f0c : data_o = 32'h44720001 ;
			32'h00100f10 : data_o = 32'h80826105 ;
			32'h00100f14 : data_o = 32'hd6227179 ;
			32'h00100f18 : data_o = 32'h87aa1800 ;
			32'h00100f1c : data_o = 32'h0fa38736 ;
			32'h00100f20 : data_o = 32'h87aefcf4 ;
			32'h00100f24 : data_o = 32'hfcf40f23 ;
			32'h00100f28 : data_o = 32'h0ea387b2 ;
			32'h00100f2c : data_o = 32'h87bafcf4 ;
			32'h00100f30 : data_o = 32'hfcf40e23 ;
			32'h00100f34 : data_o = 32'hfdf44703 ;
			32'h00100f38 : data_o = 32'hfde44783 ;
			32'h00100f3c : data_o = 32'h8f5d07a2 ;
			32'h00100f40 : data_o = 32'hfdd44783 ;
			32'h00100f44 : data_o = 32'h8f5d07c2 ;
			32'h00100f48 : data_o = 32'hfdc44783 ;
			32'h00100f4c : data_o = 32'h8fd907e2 ;
			32'h00100f50 : data_o = 32'hfef42623 ;
			32'h00100f54 : data_o = 32'h700007b7 ;
			32'h00100f58 : data_o = 32'h03478793 ;
			32'h00100f5c : data_o = 32'hfec42703 ;
			32'h00100f60 : data_o = 32'h0001c398 ;
			32'h00100f64 : data_o = 32'h61455432 ;
			32'h00100f68 : data_o = 32'h71798082 ;
			32'h00100f6c : data_o = 32'h1800d622 ;
			32'h00100f70 : data_o = 32'h873687aa ;
			32'h00100f74 : data_o = 32'hfcf40fa3 ;
			32'h00100f78 : data_o = 32'h0f2387ae ;
			32'h00100f7c : data_o = 32'h87b2fcf4 ;
			32'h00100f80 : data_o = 32'hfcf40ea3 ;
			32'h00100f84 : data_o = 32'h0e2387ba ;
			32'h00100f88 : data_o = 32'h4703fcf4 ;
			32'h00100f8c : data_o = 32'h4783fdf4 ;
			32'h00100f90 : data_o = 32'h07a2fde4 ;
			32'h00100f94 : data_o = 32'h47838f5d ;
			32'h00100f98 : data_o = 32'h07c2fdd4 ;
			32'h00100f9c : data_o = 32'h47838f5d ;
			32'h00100fa0 : data_o = 32'h07e2fdc4 ;
			32'h00100fa4 : data_o = 32'h26238fd9 ;
			32'h00100fa8 : data_o = 32'h07b7fef4 ;
			32'h00100fac : data_o = 32'h87937000 ;
			32'h00100fb0 : data_o = 32'h27030387 ;
			32'h00100fb4 : data_o = 32'hc398fec4 ;
			32'h00100fb8 : data_o = 32'h54320001 ;
			32'h00100fbc : data_o = 32'h80826145 ;
			32'h00100fc0 : data_o = 32'hce221101 ;
			32'h00100fc4 : data_o = 32'h26231000 ;
			32'h00100fc8 : data_o = 32'h07b7fea4 ;
			32'h00100fcc : data_o = 32'h87937000 ;
			32'h00100fd0 : data_o = 32'h27030207 ;
			32'h00100fd4 : data_o = 32'hc398fec4 ;
			32'h00100fd8 : data_o = 32'h44720001 ;
			32'h00100fdc : data_o = 32'h80826105 ;
			32'h00100fe0 : data_o = 32'hc6221141 ;
			32'h00100fe4 : data_o = 32'h07b70800 ;
			32'h00100fe8 : data_o = 32'h87937000 ;
			32'h00100fec : data_o = 32'h47050247 ;
			32'h00100ff0 : data_o = 32'h0001c398 ;
			32'h00100ff4 : data_o = 32'h01414432 ;
			32'h00100ff8 : data_o = 32'h11418082 ;
			32'h00100ffc : data_o = 32'h0800c622 ;
			32'h00101000 : data_o = 32'h700007b7 ;
			32'h00101004 : data_o = 32'h02878793 ;
			32'h00101008 : data_o = 32'h853e439c ;
			32'h0010100c : data_o = 32'h01414432 ;
			32'h00101010 : data_o = 32'h11418082 ;
			32'h00101014 : data_o = 32'h0800c622 ;
			32'h00101018 : data_o = 32'h700007b7 ;
			32'h0010101c : data_o = 32'h02c78793 ;
			32'h00101020 : data_o = 32'h853e439c ;
			32'h00101024 : data_o = 32'h01414432 ;
			32'h00101028 : data_o = 32'h11418082 ;
			32'h0010102c : data_o = 32'h0800c622 ;
			32'h00101030 : data_o = 32'h700007b7 ;
			32'h00101034 : data_o = 32'h03078793 ;
			32'h00101038 : data_o = 32'h853e439c ;
			32'h0010103c : data_o = 32'h01414432 ;
			32'h00101040 : data_o = 32'h11018082 ;
			32'h00101044 : data_o = 32'h1000ce22 ;
			32'h00101048 : data_o = 32'hfea42623 ;
			32'h0010104c : data_o = 32'hfec42703 ;
			32'h00101050 : data_o = 32'h700007b7 ;
			32'h00101054 : data_o = 32'h10078793 ;
			32'h00101058 : data_o = 32'h439c97ba ;
			32'h0010105c : data_o = 32'h4472853e ;
			32'h00101060 : data_o = 32'h80826105 ;
			32'h00101064 : data_o = 32'hce221101 ;
			32'h00101068 : data_o = 32'h26231000 ;
			32'h0010106c : data_o = 32'h07b7fea4 ;
			32'h00101070 : data_o = 32'h07e17000 ;
			32'h00101074 : data_o = 32'hfec42703 ;
			32'h00101078 : data_o = 32'h0001c398 ;
			32'h0010107c : data_o = 32'h61054472 ;
			32'h00101080 : data_o = 32'h11018082 ;
			32'h00101084 : data_o = 32'h1000ce22 ;
			32'h00101088 : data_o = 32'hfea42623 ;
			32'h0010108c : data_o = 32'h700007b7 ;
			32'h00101090 : data_o = 32'h03c78793 ;
			32'h00101094 : data_o = 32'hfec42703 ;
			32'h00101098 : data_o = 32'h0001c398 ;
			32'h0010109c : data_o = 32'h61054472 ;
			32'h001010a0 : data_o = 32'h11018082 ;
			32'h001010a4 : data_o = 32'h1000ce22 ;
			32'h001010a8 : data_o = 32'hfea42623 ;
			32'h001010ac : data_o = 32'h873687ae ;
			32'h001010b0 : data_o = 32'hfef405a3 ;
			32'h001010b4 : data_o = 32'h052387b2 ;
			32'h001010b8 : data_o = 32'h87bafef4 ;
			32'h001010bc : data_o = 32'hfef404a3 ;
			32'h001010c0 : data_o = 32'hfeb44783 ;
			32'h001010c4 : data_o = 32'hf713078e ;
			32'h001010c8 : data_o = 32'h47830187 ;
			32'h001010cc : data_o = 32'h0796fea4 ;
			32'h001010d0 : data_o = 32'h47838f5d ;
			32'h001010d4 : data_o = 32'h078afe94 ;
			32'h001010d8 : data_o = 32'h8f5d8b91 ;
			32'h001010dc : data_o = 32'h700007b7 ;
			32'h001010e0 : data_o = 32'h10078793 ;
			32'h001010e4 : data_o = 32'h873e97ba ;
			32'h001010e8 : data_o = 32'hfec42783 ;
			32'h001010ec : data_o = 32'hfff7c793 ;
			32'h001010f0 : data_o = 32'h0001c31c ;
			32'h001010f4 : data_o = 32'h61054472 ;
			32'h001010f8 : data_o = 32'hf06f8082 ;
			32'h001010fc : data_o = 32'h0093a2ff ;
			32'h00101100 : data_o = 32'h81060000 ;
			32'h00101104 : data_o = 32'h82068186 ;
			32'h00101108 : data_o = 32'h83068286 ;
			32'h0010110c : data_o = 32'h84068386 ;
			32'h00101110 : data_o = 32'h85068486 ;
			32'h00101114 : data_o = 32'h86068586 ;
			32'h00101118 : data_o = 32'h87068686 ;
			32'h0010111c : data_o = 32'h88068786 ;
			32'h00101120 : data_o = 32'h89068886 ;
			32'h00101124 : data_o = 32'h8a068986 ;
			32'h00101128 : data_o = 32'h8b068a86 ;
			32'h0010112c : data_o = 32'h8c068b86 ;
			32'h00101130 : data_o = 32'h8d068c86 ;
			32'h00101134 : data_o = 32'h8e068d86 ;
			32'h00101138 : data_o = 32'h8f068e86 ;
			32'h0010113c : data_o = 32'hf1178f86 ;
			32'h00101140 : data_o = 32'h01130011 ;
			32'h00101144 : data_o = 32'hfd17ec21 ;
			32'h00101148 : data_o = 32'h0d13000f ;
			32'h0010114c : data_o = 32'hfd97ec2d ;
			32'h00101150 : data_o = 32'h8d93000f ;
			32'h00101154 : data_o = 32'h5763ee2d ;
			32'h00101158 : data_o = 32'h202301bd ;
			32'h0010115c : data_o = 32'h0d11000d ;
			32'h00101160 : data_o = 32'hffaddde3 ;
			32'h00101164 : data_o = 32'h45814501 ;
			32'h00101168 : data_o = 32'ha66ff0ef ;
			32'h0010116c : data_o = 32'h000202b7 ;
			32'h00101170 : data_o = 32'h430502a1 ;
			32'h00101174 : data_o = 32'h0062a023 ;
			32'h00101178 : data_o = 32'h10500073 ;
			32'h0010117c : data_o = 32'h47b3bff5 ;
			32'h00101180 : data_o = 32'h8b8d00b5 ;
			32'h00101184 : data_o = 32'h00c508b3 ;
			32'h00101188 : data_o = 32'h478de7b1 ;
			32'h0010118c : data_o = 32'h04c7f463 ;
			32'h00101190 : data_o = 32'h00357793 ;
			32'h00101194 : data_o = 32'hebb9872a ;
			32'h00101198 : data_o = 32'hffc8f613 ;
			32'h0010119c : data_o = 32'h40e606b3 ;
			32'h001011a0 : data_o = 32'h02000793 ;
			32'h001011a4 : data_o = 32'h06d7c863 ;
			32'h001011a8 : data_o = 32'h87ba86ae ;
			32'h001011ac : data_o = 32'h02c77163 ;
			32'h001011b0 : data_o = 32'h0006a803 ;
			32'h001011b4 : data_o = 32'h06910791 ;
			32'h001011b8 : data_o = 32'hff07ae23 ;
			32'h001011bc : data_o = 32'hfec7eae3 ;
			32'h001011c0 : data_o = 32'hfff60793 ;
			32'h001011c4 : data_o = 32'h9bf18f99 ;
			32'h001011c8 : data_o = 32'h973e0791 ;
			32'h001011cc : data_o = 32'h666395be ;
			32'h001011d0 : data_o = 32'h80820117 ;
			32'h001011d4 : data_o = 32'h7e63872a ;
			32'h001011d8 : data_o = 32'hc7830315 ;
			32'h001011dc : data_o = 32'h07050005 ;
			32'h001011e0 : data_o = 32'h0fa30585 ;
			32'h001011e4 : data_o = 32'h9ae3fef7 ;
			32'h001011e8 : data_o = 32'h8082fee8 ;
			32'h001011ec : data_o = 32'h0005c683 ;
			32'h001011f0 : data_o = 32'h77930705 ;
			32'h001011f4 : data_o = 32'h0fa30037 ;
			32'h001011f8 : data_o = 32'h0585fed7 ;
			32'h001011fc : data_o = 32'hc683dfd1 ;
			32'h00101200 : data_o = 32'h07050005 ;
			32'h00101204 : data_o = 32'h00377793 ;
			32'h00101208 : data_o = 32'hfed70fa3 ;
			32'h0010120c : data_o = 32'hfff90585 ;
			32'h00101210 : data_o = 32'h8082b761 ;
			32'h00101214 : data_o = 32'hc6221141 ;
			32'h00101218 : data_o = 32'h02000413 ;
			32'h0010121c : data_o = 32'h0005a383 ;
			32'h00101220 : data_o = 32'h0045a283 ;
			32'h00101224 : data_o = 32'h0085af83 ;
			32'h00101228 : data_o = 32'h00c5af03 ;
			32'h0010122c : data_o = 32'h0105ae83 ;
			32'h00101230 : data_o = 32'h0145ae03 ;
			32'h00101234 : data_o = 32'h0185a303 ;
			32'h00101238 : data_o = 32'h01c5a803 ;
			32'h0010123c : data_o = 32'h07135194 ;
			32'h00101240 : data_o = 32'h07b30247 ;
			32'h00101244 : data_o = 32'h2e2340e6 ;
			32'h00101248 : data_o = 32'h2023fc77 ;
			32'h0010124c : data_o = 32'h2223fe57 ;
			32'h00101250 : data_o = 32'h2423fff7 ;
			32'h00101254 : data_o = 32'h2623ffe7 ;
			32'h00101258 : data_o = 32'h2823ffd7 ;
			32'h0010125c : data_o = 32'h2a23ffc7 ;
			32'h00101260 : data_o = 32'h2c23fe67 ;
			32'h00101264 : data_o = 32'h2e23ff07 ;
			32'h00101268 : data_o = 32'h8593fed7 ;
			32'h0010126c : data_o = 32'h47e30245 ;
			32'h00101270 : data_o = 32'h86aefaf4 ;
			32'h00101274 : data_o = 32'h716387ba ;
			32'h00101278 : data_o = 32'ha80302c7 ;
			32'h0010127c : data_o = 32'h07910006 ;
			32'h00101280 : data_o = 32'hae230691 ;
			32'h00101284 : data_o = 32'heae3ff07 ;
			32'h00101288 : data_o = 32'h0793fec7 ;
			32'h0010128c : data_o = 32'h8f99fff6 ;
			32'h00101290 : data_o = 32'h07919bf1 ;
			32'h00101294 : data_o = 32'h95be973e ;
			32'h00101298 : data_o = 32'h01176563 ;
			32'h0010129c : data_o = 32'h01414432 ;
			32'h001012a0 : data_o = 32'hc7838082 ;
			32'h001012a4 : data_o = 32'h07050005 ;
			32'h001012a8 : data_o = 32'h0fa30585 ;
			32'h001012ac : data_o = 32'h87e3fef7 ;
			32'h001012b0 : data_o = 32'hc783fee8 ;
			32'h001012b4 : data_o = 32'h07050005 ;
			32'h001012b8 : data_o = 32'h0fa30585 ;
			32'h001012bc : data_o = 32'h92e3fef7 ;
			32'h001012c0 : data_o = 32'hbfe9fee8 ;
			32'h001012c4 : data_o = 32'h50505553 ;
			32'h001012c8 : data_o = 32'h465f594c ;
			32'h001012cc : data_o = 32'h0a4d524f ;
			32'h001012d0 : data_o = 32'h00000000 ;
			32'h001012d4 : data_o = 32'h50505553 ;
			32'h001012d8 : data_o = 32'h535f594c ;
			32'h001012dc : data_o = 32'h000a5445 ;
			32'h001012e0 : data_o = 32'h50505553 ;
			32'h001012e4 : data_o = 32'h525f594c ;
			32'h001012e8 : data_o = 32'h54455345 ;
			32'h001012ec : data_o = 32'h0000000a ;
			32'h001012f0 : data_o = 32'h50505553 ;
			32'h001012f4 : data_o = 32'h525f594c ;
			32'h001012f8 : data_o = 32'h0a444145 ;
			32'h001012fc : data_o = 32'h00000000 ;
			32'h00101300 : data_o = 32'h52415453 ;
			32'h00101304 : data_o = 32'h52415f54 ;
			32'h00101308 : data_o = 32'h0a594152 ;
			32'h0010130c : data_o = 32'h00000000 ;
			32'h00101310 : data_o = 32'h5f444e45 ;
			32'h00101314 : data_o = 32'h41525241 ;
			32'h00101318 : data_o = 32'h00000a59 ;
			32'h0010131c : data_o = 32'h0a444e45 ;
			32'h00101320 : data_o = 32'h00000000 ;
			32'h00101324 : data_o = 32'h00000000 ;
			32'h00101328 : data_o = 32'h00000000 ;
			32'h0010132c : data_o = 32'h00000000 ;
			32'h00101330 : data_o = 32'h00000000 ;
			32'h00101334 : data_o = 32'h00000000 ;
			32'h00101338 : data_o = 32'h00000000 ;
			32'h0010133c : data_o = 32'h00000000 ;
			32'h00101340 : data_o = 32'h00000000 ;
			32'h00101344 : data_o = 32'h00000000 ;
			32'h00101348 : data_o = 32'h00000000 ;
			32'h0010134c : data_o = 32'h00000000 ;
			32'h00101350 : data_o = 32'h00000000 ;
			32'h00101354 : data_o = 32'h00000000 ;
			32'h00101358 : data_o = 32'h00000000 ;
			32'h0010135c : data_o = 32'hff070000 ;
			32'h00101360 : data_o = 32'h0000e0ff ;
			32'h00101364 : data_o = 32'hff070000 ;
			32'h00101368 : data_o = 32'h0000e0ff ;
			32'h0010136c : data_o = 32'hff070000 ;
			32'h00101370 : data_o = 32'h0000e0ff ;
			32'h00101374 : data_o = 32'hff070000 ;
			32'h00101378 : data_o = 32'h0000e0ff ;
			32'h0010137c : data_o = 32'hffff0300 ;
			32'h00101380 : data_o = 32'h00c0ffff ;
			32'h00101384 : data_o = 32'hffff0300 ;
			32'h00101388 : data_o = 32'h00c0ffff ;
			32'h0010138c : data_o = 32'hffff0300 ;
			32'h00101390 : data_o = 32'h00c0ffff ;
			32'h00101394 : data_o = 32'hffc71f00 ;
			32'h00101398 : data_o = 32'h00f8e3ff ;
			32'h0010139c : data_o = 32'hffc71f00 ;
			32'h001013a0 : data_o = 32'h00f8e3ff ;
			32'h001013a4 : data_o = 32'hffc71f00 ;
			32'h001013a8 : data_o = 32'h00f8e3ff ;
			32'h001013ac : data_o = 32'hffc71f00 ;
			32'h001013b0 : data_o = 32'h00f8e3ff ;
			32'h001013b4 : data_o = 32'hffc7ff01 ;
			32'h001013b8 : data_o = 32'h80ffe3ff ;
			32'h001013bc : data_o = 32'hffc7ff01 ;
			32'h001013c0 : data_o = 32'h80ffe3ff ;
			32'h001013c4 : data_o = 32'hffc7ff01 ;
			32'h001013c8 : data_o = 32'h80ffe3ff ;
			32'h001013cc : data_o = 32'hffc7ff01 ;
			32'h001013d0 : data_o = 32'h80ffe3ff ;
			32'h001013d4 : data_o = 32'hffc7ff01 ;
			32'h001013d8 : data_o = 32'h80ffe3ff ;
			32'h001013dc : data_o = 32'hffc7ff01 ;
			32'h001013e0 : data_o = 32'h80ffe3ff ;
			32'h001013e4 : data_o = 32'hffc7ff01 ;
			32'h001013e8 : data_o = 32'h80ffe3ff ;
			32'h001013ec : data_o = 32'h7ff8ff0f ;
			32'h001013f0 : data_o = 32'hf0ff1ffe ;
			32'h001013f4 : data_o = 32'h7ff8ff0f ;
			32'h001013f8 : data_o = 32'hf0ff1ffe ;
			32'h001013fc : data_o = 32'h7ff8ff0f ;
			32'h00101400 : data_o = 32'hf0ff1ffe ;
			32'h00101404 : data_o = 32'h00f81f0e ;
			32'h00101408 : data_o = 32'h70f81f00 ;
			32'h0010140c : data_o = 32'h00f81f0e ;
			32'h00101410 : data_o = 32'h70f81f00 ;
			32'h00101414 : data_o = 32'h00f81f0e ;
			32'h00101418 : data_o = 32'h70f81f00 ;
			32'h0010141c : data_o = 32'h00f81f0e ;
			32'h00101420 : data_o = 32'h70f81f00 ;
			32'h00101424 : data_o = 32'h0000e00f ;
			32'h00101428 : data_o = 32'hf0070000 ;
			32'h0010142c : data_o = 32'h0000e00f ;
			32'h00101430 : data_o = 32'hf0070000 ;
			32'h00101434 : data_o = 32'h0000e00f ;
			32'h00101438 : data_o = 32'hf0070000 ;
			32'h0010143c : data_o = 32'h0000e00f ;
			32'h00101440 : data_o = 32'hf0070000 ;
			32'h00101444 : data_o = 32'h7f00e00f ;
			32'h00101448 : data_o = 32'hf00700fe ;
			32'h0010144c : data_o = 32'h7f00e00f ;
			32'h00101450 : data_o = 32'hf00700fe ;
			32'h00101454 : data_o = 32'h7f00e00f ;
			32'h00101458 : data_o = 32'hf00700fe ;
			32'h0010145c : data_o = 32'h8007fc0f ;
			32'h00101460 : data_o = 32'hf03fe001 ;
			32'h00101464 : data_o = 32'h8007fc0f ;
			32'h00101468 : data_o = 32'hf03fe001 ;
			32'h0010146c : data_o = 32'h8007fc0f ;
			32'h00101470 : data_o = 32'hf03fe001 ;
			32'h00101474 : data_o = 32'h8007fc0f ;
			32'h00101478 : data_o = 32'hf03fe001 ;
			32'h0010147c : data_o = 32'h0038fc0f ;
			32'h00101480 : data_o = 32'hf03f1c00 ;
			32'h00101484 : data_o = 32'h0038fc0f ;
			32'h00101488 : data_o = 32'hf03f1c00 ;
			32'h0010148c : data_o = 32'h0038fc0f ;
			32'h00101490 : data_o = 32'hf03f1c00 ;
			32'h00101494 : data_o = 32'h00f8e30f ;
			32'h00101498 : data_o = 32'hf0c71f00 ;
			32'h0010149c : data_o = 32'h00f8e30f ;
			32'h001014a0 : data_o = 32'hf0c71f00 ;
			32'h001014a4 : data_o = 32'h00f8e30f ;
			32'h001014a8 : data_o = 32'hf0c71f00 ;
			32'h001014ac : data_o = 32'h00f8e30f ;
			32'h001014b0 : data_o = 32'hf0c71f00 ;
			32'h001014b4 : data_o = 32'h00c0ff01 ;
			32'h001014b8 : data_o = 32'h80ff0300 ;
			32'h001014bc : data_o = 32'h00c0ff01 ;
			32'h001014c0 : data_o = 32'h80ff0300 ;
			32'h001014c4 : data_o = 32'h00c0ff01 ;
			32'h001014c8 : data_o = 32'h80ff0300 ;
			32'h001014cc : data_o = 32'h00000000 ;
			32'h001014d0 : data_o = 32'h00000000 ;
			32'h001014d4 : data_o = 32'h00000000 ;
			32'h001014d8 : data_o = 32'h00000000 ;
			32'h001014dc : data_o = 32'h00000000 ;
			32'h001014e0 : data_o = 32'h00000000 ;
			32'h001014e4 : data_o = 32'h00000000 ;
			32'h001014e8 : data_o = 32'h00000000 ;
			32'h001014ec : data_o = 32'h00000000 ;
			32'h001014f0 : data_o = 32'h00000000 ;
			32'h001014f4 : data_o = 32'h00000000 ;
			32'h001014f8 : data_o = 32'h00000000 ;
			32'h001014fc : data_o = 32'h00000000 ;
			32'h00101500 : data_o = 32'h00000000 ;
			32'h00101504 : data_o = 32'h00000000 ;
			32'h00101508 : data_o = 32'h00000000 ;
			32'h0010150c : data_o = 32'h00000000 ;
			32'h00101510 : data_o = 32'h00000000 ;
			32'h00101514 : data_o = 32'h00000000 ;
			32'h00101518 : data_o = 32'h00000000 ;
			32'h0010151c : data_o = 32'h00000000 ;
			32'h00101520 : data_o = 32'h00000000 ;
			32'h00101524 : data_o = 32'h45435845 ;
			32'h00101528 : data_o = 32'h4f495450 ;
			32'h0010152c : data_o = 32'h2121214e ;
			32'h00101530 : data_o = 32'h0000000a ;
			32'h00101534 : data_o = 32'h3d3d3d3d ;
			32'h00101538 : data_o = 32'h3d3d3d3d ;
			32'h0010153c : data_o = 32'h3d3d3d3d ;
			32'h00101540 : data_o = 32'h0000000a ;
			32'h00101544 : data_o = 32'h4350454d ;
			32'h00101548 : data_o = 32'h2020203a ;
			32'h0010154c : data_o = 32'h00007830 ;
			32'h00101550 : data_o = 32'h41434d0a ;
			32'h00101554 : data_o = 32'h3a455355 ;
			32'h00101558 : data_o = 32'h00783020 ;
			32'h0010155c : data_o = 32'h56544d0a ;
			32'h00101560 : data_o = 32'h203a4c41 ;
			32'h00101564 : data_o = 32'h00783020 ;
			32'h00101568 : data_o = 32'h00100000 ;
			default : data_o = 32'h00000000 ;
		endcase 
	end
endmodule
